
module mux_top ( out, in1, in2, sel );
  input in1, in2, sel;
  output out;
  wire   n2, n3, n4;

  AND2XLTH U4 ( .A(in1), .B(sel), .Y(n2) );
  OR2XLTH U2 ( .A(n2), .B(n3), .Y(out) );
  AND2XLTH U3 ( .A(in2), .B(n4), .Y(n3) );
  INVXLTH U1 ( .A(sel), .Y(n4) );
endmodule


module counter_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXLTH U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXLTH U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXLTH U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXLTH U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXLTH U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR2XLTH U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVXLTH U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module counter_test_1 ( out1, sel, clk, rst, test_si, test_so, test_se );
  input [1:0] sel;
  input clk, rst, test_si, test_se;
  output out1, test_so;
  wire   N18, N19, N20, N21, N22, N23, N24, n25, n26, n27, n28, n29, n30, n31,
         n32, n9, n10, n6, n7, n8, n11, n12, n13, n14, n15, n42, n43, n44, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58;
  wire   [6:0] count;

  counter_DW01_inc_0 r310 ( .A({count[6], n55, count[4:2], n57, count[0]}), 
        .SUM({N24, N23, N22, N21, N20, N19, N18}) );
  SDFFRQXLTH count_reg_1_ ( .D(n26), .SI(count[0]), .SE(n52), .CK(clk), .RN(
        rst), .Q(count[1]) );
  SDFFRQX1TH count_reg_0_ ( .D(n32), .SI(test_si), .SE(n52), .CK(clk), .RN(rst), .Q(count[0]) );
  SDFFRQX1TH count_reg_2_ ( .D(n27), .SI(n57), .SE(n53), .CK(clk), .RN(rst), 
        .Q(count[2]) );
  SDFFRQX1TH count_reg_5_ ( .D(n30), .SI(count[4]), .SE(n50), .CK(clk), .RN(
        rst), .Q(count[5]) );
  SDFFRQX1TH count_reg_6_ ( .D(n31), .SI(n55), .SE(n51), .CK(clk), .RN(rst), 
        .Q(count[6]) );
  SDFFSRXLTH out1_reg ( .D(n25), .SI(n54), .SE(n53), .CK(clk), .SN(1'b1), .RN(
        rst), .Q(out1), .QN(test_so) );
  SDFFRX1TH count_reg_3_ ( .D(n28), .SI(count[2]), .SE(n50), .CK(clk), .RN(rst), .Q(count[3]), .QN(n9) );
  SDFFRX1TH count_reg_4_ ( .D(n29), .SI(count[3]), .SE(n51), .CK(clk), .RN(rst), .Q(count[4]), .QN(n10) );
  NAND2XLTH U5 ( .A(n13), .B(n44), .Y(n12) );
  INVXLTH U6 ( .A(count[5]), .Y(n44) );
  INVXLTH U7 ( .A(count[2]), .Y(n43) );
  OAI21X6TH U8 ( .A0(sel[1]), .A1(n7), .B0(n8), .Y(n6) );
  AOI211X1TH U9 ( .A0(n14), .A1(count[5]), .B0(count[6]), .C0(n15), .Y(n7) );
  NOR3XLTH U10 ( .A(n10), .B(sel[0]), .C(n9), .Y(n11) );
  CLKINVX2TH U11 ( .A(n6), .Y(n42) );
  AO22XLTH U12 ( .A0(n54), .A1(n6), .B0(N24), .B1(n42), .Y(n31) );
  AO22XLTH U13 ( .A0(count[0]), .A1(n6), .B0(N18), .B1(n42), .Y(n32) );
  OR2XLTH U14 ( .A(out1), .B(n6), .Y(n25) );
  AO22XLTH U15 ( .A0(n58), .A1(n6), .B0(N19), .B1(n42), .Y(n26) );
  AOI211XLTH U16 ( .A0(n9), .A1(n43), .B0(sel[0]), .C0(n10), .Y(n15) );
  NAND2XLTH U17 ( .A(n9), .B(n13), .Y(n14) );
  OAI2B2XLTH U18 ( .A1N(N23), .A0(n6), .B0(n42), .B1(n44), .Y(n30) );
  OAI2B2XLTH U19 ( .A1N(N20), .A0(n6), .B0(n42), .B1(n43), .Y(n27) );
  AOI32XLTH U20 ( .A0(count[5]), .A1(count[2]), .A2(n11), .B0(count[6]), .B1(
        n12), .Y(n8) );
  OAI2B2XLTH U21 ( .A1N(N21), .A0(n6), .B0(n9), .B1(n42), .Y(n28) );
  OAI2B2XLTH U22 ( .A1N(N22), .A0(n6), .B0(n10), .B1(n42), .Y(n29) );
  AND2XLTH U23 ( .A(sel[0]), .B(n10), .Y(n13) );
  INVXLTH U39 ( .A(test_se), .Y(n48) );
  INVXLTH U40 ( .A(test_se), .Y(n49) );
  INVXLTH U41 ( .A(n48), .Y(n50) );
  INVXLTH U42 ( .A(n48), .Y(n51) );
  INVXLTH U43 ( .A(n49), .Y(n52) );
  INVXLTH U44 ( .A(n49), .Y(n53) );
  DLY1X1TH U45 ( .A(count[6]), .Y(n54) );
  DLY1X1TH U46 ( .A(count[5]), .Y(n55) );
  INVXLTH U47 ( .A(count[1]), .Y(n56) );
  INVXLTH U48 ( .A(n56), .Y(n57) );
  INVXLTH U49 ( .A(n56), .Y(n58) );
endmodule


module counter_PISO_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  ADDHXLTH U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXLTH U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXLTH U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXLTH U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXLTH U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXLTH U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXLTH U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXLTH U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVXLTH U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2XLTH U2 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
endmodule


module counter_PISO_DW01_inc_1 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  ADDHXLTH U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXLTH U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXLTH U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXLTH U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXLTH U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXLTH U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXLTH U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXLTH U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  INVXLTH U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2XLTH U2 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
endmodule


module mux1_test_0 ( out, in1, in2, sel, clk, rst, test_si, test_se );
  input in1, in2, sel, clk, rst, test_si, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(test_si), .SE(test_se), .CK(clk), .RN(rst), 
        .Q(out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_1 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_2 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_3 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_4 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_5 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_6 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_7 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_8 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_9 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_10 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_11 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_12 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_13 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_14 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_15 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_16 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_17 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_18 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_19 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_20 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_21 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_22 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_23 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_24 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_25 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_26 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_27 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_28 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_29 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_30 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_31 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_32 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_33 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_34 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_35 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_36 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_37 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_38 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_39 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_40 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_41 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_42 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_43 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_44 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_45 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_46 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module mux1_test_47 ( out, in1, in2, sel, clk, rst, test_se );
  input in1, in2, sel, clk, rst, test_se;
  output out;
  wire   N2;

  SDFFRQXLTH out_reg ( .D(N2), .SI(in1), .SE(test_se), .CK(clk), .RN(rst), .Q(
        out) );
  AO2B2XLTH U3 ( .B0(sel), .B1(in1), .A0(in2), .A1N(sel), .Y(N2) );
endmodule


module PISO_test_1 ( out, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, 
        in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, 
        in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, 
        in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, 
        in47, in48, sel, clk, rst, test_si, test_so, test_se );
  input in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13,
         in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24,
         in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35,
         in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46,
         in47, in48, sel, clk, rst, test_si, test_se;
  output out, test_so;
  wire   t1, t2, t3, t4, t5, t6, t7, t8, t9, t10, t11, t12, t13, t14, t15, t16,
         t17, t18, t19, t20, t21, t22, t23, t24, t25, t26, t27, t28, t29, t30,
         t31, t32, t33, t34, t35, t36, t37, t38, t39, t40, t41, t42, t43, t44,
         t45, t46, t47, t48, n13, n14, n15, n16, n17, n18, n19, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55;

  mux1_test_0 mux1_1 ( .out(t1), .in1(in48), .in2(in48), .sel(n19), .clk(clk), 
        .rst(n16), .test_si(test_si), .test_se(n50) );
  mux1_test_1 mux1_2 ( .out(t2), .in1(t1), .in2(in47), .sel(n17), .clk(clk), 
        .rst(n13), .test_se(n50) );
  mux1_test_2 mux1_3 ( .out(t3), .in1(t2), .in2(in46), .sel(n17), .clk(clk), 
        .rst(n13), .test_se(n49) );
  mux1_test_3 mux1_4 ( .out(t4), .in1(t3), .in2(in45), .sel(n17), .clk(clk), 
        .rst(n13), .test_se(n50) );
  mux1_test_4 mux1_5 ( .out(t5), .in1(t4), .in2(in44), .sel(n17), .clk(clk), 
        .rst(n13), .test_se(n49) );
  mux1_test_5 mux1_6 ( .out(t6), .in1(t5), .in2(in43), .sel(n17), .clk(clk), 
        .rst(n13), .test_se(n49) );
  mux1_test_6 mux1_7 ( .out(t7), .in1(t6), .in2(in42), .sel(n17), .clk(clk), 
        .rst(n13), .test_se(n48) );
  mux1_test_7 mux1_8 ( .out(t8), .in1(t7), .in2(in41), .sel(n17), .clk(clk), 
        .rst(n13), .test_se(n49) );
  mux1_test_8 mux1_9 ( .out(t9), .in1(t8), .in2(in40), .sel(n17), .clk(clk), 
        .rst(n13), .test_se(n48) );
  mux1_test_9 mux1_10 ( .out(t10), .in1(t9), .in2(in39), .sel(n17), .clk(clk), 
        .rst(n13), .test_se(n48) );
  mux1_test_10 mux1_11 ( .out(t11), .in1(t10), .in2(in38), .sel(n17), .clk(clk), .rst(n13), .test_se(n45) );
  mux1_test_11 mux1_12 ( .out(t12), .in1(t11), .in2(in37), .sel(n17), .clk(clk), .rst(n13), .test_se(n48) );
  mux1_test_12 mux1_13 ( .out(t13), .in1(t12), .in2(in36), .sel(n17), .clk(clk), .rst(n13), .test_se(n45) );
  mux1_test_13 mux1_14 ( .out(t14), .in1(t13), .in2(in35), .sel(n17), .clk(clk), .rst(n14), .test_se(n45) );
  mux1_test_14 mux1_15 ( .out(t15), .in1(t14), .in2(in34), .sel(n18), .clk(clk), .rst(n14), .test_se(n46) );
  mux1_test_15 mux1_16 ( .out(t16), .in1(t15), .in2(in33), .sel(n18), .clk(clk), .rst(n14), .test_se(n45) );
  mux1_test_16 mux1_17 ( .out(t17), .in1(t16), .in2(in32), .sel(n18), .clk(clk), .rst(n14), .test_se(n46) );
  mux1_test_17 mux1_18 ( .out(t18), .in1(t17), .in2(in31), .sel(n18), .clk(clk), .rst(n14), .test_se(n46) );
  mux1_test_18 mux1_19 ( .out(t19), .in1(t18), .in2(in30), .sel(n18), .clk(clk), .rst(n14), .test_se(n47) );
  mux1_test_19 mux1_20 ( .out(t20), .in1(t19), .in2(in29), .sel(n18), .clk(clk), .rst(n14), .test_se(n46) );
  mux1_test_20 mux1_21 ( .out(t21), .in1(t20), .in2(in28), .sel(n18), .clk(clk), .rst(n14), .test_se(n47) );
  mux1_test_21 mux1_22 ( .out(t22), .in1(t21), .in2(in27), .sel(n18), .clk(clk), .rst(n14), .test_se(n47) );
  mux1_test_22 mux1_23 ( .out(t23), .in1(t22), .in2(in26), .sel(n18), .clk(clk), .rst(n14), .test_se(n26) );
  mux1_test_23 mux1_24 ( .out(t24), .in1(t23), .in2(in25), .sel(n18), .clk(clk), .rst(n14), .test_se(n27) );
  mux1_test_24 mux1_25 ( .out(t25), .in1(t24), .in2(in24), .sel(n18), .clk(clk), .rst(n14), .test_se(n28) );
  mux1_test_25 mux1_26 ( .out(t26), .in1(t25), .in2(in23), .sel(n18), .clk(clk), .rst(n15), .test_se(n25) );
  mux1_test_26 mux1_27 ( .out(t27), .in1(t26), .in2(in22), .sel(n18), .clk(clk), .rst(n15), .test_se(n26) );
  mux1_test_27 mux1_28 ( .out(t28), .in1(t27), .in2(in21), .sel(n19), .clk(clk), .rst(n15), .test_se(n30) );
  mux1_test_28 mux1_29 ( .out(t29), .in1(t28), .in2(in20), .sel(n19), .clk(clk), .rst(n15), .test_se(n31) );
  mux1_test_29 mux1_30 ( .out(t30), .in1(t29), .in2(in19), .sel(n19), .clk(clk), .rst(n15), .test_se(n32) );
  mux1_test_30 mux1_31 ( .out(t31), .in1(t30), .in2(in18), .sel(n19), .clk(clk), .rst(n15), .test_se(n29) );
  mux1_test_31 mux1_32 ( .out(t32), .in1(t31), .in2(in17), .sel(n19), .clk(clk), .rst(n15), .test_se(n30) );
  mux1_test_32 mux1_33 ( .out(t33), .in1(t32), .in2(in16), .sel(n19), .clk(clk), .rst(n15), .test_se(n34) );
  mux1_test_33 mux1_34 ( .out(t34), .in1(t33), .in2(in15), .sel(n19), .clk(clk), .rst(n15), .test_se(n35) );
  mux1_test_34 mux1_35 ( .out(t35), .in1(t34), .in2(in14), .sel(n19), .clk(clk), .rst(n15), .test_se(n36) );
  mux1_test_35 mux1_36 ( .out(t36), .in1(t35), .in2(in13), .sel(n19), .clk(clk), .rst(n15), .test_se(n33) );
  mux1_test_36 mux1_37 ( .out(t37), .in1(t36), .in2(in12), .sel(n19), .clk(clk), .rst(n15), .test_se(n34) );
  mux1_test_37 mux1_38 ( .out(t38), .in1(t37), .in2(in11), .sel(n19), .clk(clk), .rst(n16), .test_se(n38) );
  mux1_test_38 mux1_39 ( .out(t39), .in1(t38), .in2(in10), .sel(n19), .clk(clk), .rst(n16), .test_se(n39) );
  mux1_test_39 mux1_40 ( .out(t40), .in1(t39), .in2(in9), .sel(n19), .clk(clk), 
        .rst(n16), .test_se(n40) );
  mux1_test_40 mux1_41 ( .out(t41), .in1(t40), .in2(in8), .sel(n17), .clk(clk), 
        .rst(n16), .test_se(n37) );
  mux1_test_41 mux1_42 ( .out(t42), .in1(t41), .in2(in7), .sel(n18), .clk(clk), 
        .rst(n16), .test_se(n38) );
  mux1_test_42 mux1_43 ( .out(t43), .in1(t42), .in2(in6), .sel(n18), .clk(clk), 
        .rst(n16), .test_se(n41) );
  mux1_test_43 mux1_44 ( .out(t44), .in1(t43), .in2(in5), .sel(n17), .clk(clk), 
        .rst(n16), .test_se(n42) );
  mux1_test_44 mux1_45 ( .out(t45), .in1(t44), .in2(in4), .sel(n19), .clk(clk), 
        .rst(n16), .test_se(n43) );
  mux1_test_45 mux1_46 ( .out(t46), .in1(t45), .in2(in3), .sel(n19), .clk(clk), 
        .rst(n16), .test_se(n44) );
  mux1_test_46 mux1_47 ( .out(t47), .in1(t46), .in2(in2), .sel(n19), .clk(clk), 
        .rst(n16), .test_se(n41) );
  mux1_test_47 mux1_48 ( .out(t48), .in1(t47), .in2(in1), .sel(n19), .clk(clk), 
        .rst(n16), .test_se(n42) );
  SDFFTRXLTH out_reg ( .RN(rst), .D(t48), .SI(t48), .SE(n47), .CK(clk), .Q(out), .QN(test_so) );
  CLKBUFX8TH U4 ( .A(sel), .Y(n17) );
  CLKBUFX8TH U5 ( .A(sel), .Y(n18) );
  CLKBUFX8TH U6 ( .A(sel), .Y(n19) );
  BUFX3TH U7 ( .A(rst), .Y(n13) );
  BUFX3TH U8 ( .A(rst), .Y(n14) );
  BUFX3TH U9 ( .A(rst), .Y(n15) );
  BUFX3TH U10 ( .A(rst), .Y(n16) );
  DLY1X1TH U12 ( .A(test_se), .Y(n24) );
  DLY1X1TH U13 ( .A(n51), .Y(n25) );
  DLY1X1TH U14 ( .A(n51), .Y(n26) );
  DLY1X1TH U15 ( .A(n51), .Y(n27) );
  DLY1X1TH U16 ( .A(n51), .Y(n28) );
  DLY1X1TH U17 ( .A(n52), .Y(n29) );
  DLY1X1TH U18 ( .A(n52), .Y(n30) );
  DLY1X1TH U19 ( .A(n52), .Y(n31) );
  DLY1X1TH U20 ( .A(n52), .Y(n32) );
  DLY1X1TH U21 ( .A(n53), .Y(n33) );
  DLY1X1TH U22 ( .A(n53), .Y(n34) );
  DLY1X1TH U23 ( .A(n53), .Y(n35) );
  DLY1X1TH U24 ( .A(n53), .Y(n36) );
  DLY1X1TH U25 ( .A(n54), .Y(n37) );
  DLY1X1TH U26 ( .A(n54), .Y(n38) );
  DLY1X1TH U27 ( .A(n54), .Y(n39) );
  DLY1X1TH U28 ( .A(n54), .Y(n40) );
  DLY1X1TH U29 ( .A(n55), .Y(n41) );
  DLY1X1TH U30 ( .A(n55), .Y(n42) );
  DLY1X1TH U31 ( .A(n55), .Y(n43) );
  DLY1X1TH U32 ( .A(n55), .Y(n44) );
  DLY1X1TH U33 ( .A(test_se), .Y(n45) );
  DLY1X1TH U34 ( .A(test_se), .Y(n46) );
  DLY1X1TH U35 ( .A(n24), .Y(n47) );
  DLY1X1TH U36 ( .A(n24), .Y(n48) );
  DLY1X1TH U37 ( .A(n24), .Y(n49) );
  DLY1X1TH U38 ( .A(test_se), .Y(n50) );
  DLY1X1TH U39 ( .A(n50), .Y(n51) );
  DLY1X1TH U40 ( .A(n25), .Y(n52) );
  DLY1X1TH U41 ( .A(n29), .Y(n53) );
  DLY1X1TH U42 ( .A(n33), .Y(n54) );
  DLY1X1TH U43 ( .A(n37), .Y(n55) );
endmodule


module counter_PISO_test_1 ( error, counter, hd_end, out1, in1, in2, in3, in4, 
        in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, 
        in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, 
        in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, 
        in41, in42, in43, in44, in45, in46, in47, in48, rst, ex_clk, w3, 
        test_si, test_se );
  output [9:0] error;
  output [9:0] counter;
  input in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13,
         in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24,
         in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35,
         in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46,
         in47, in48, rst, ex_clk, w3, test_si, test_se;
  output hd_end, out1;
  wire   w2, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N18, N19, N20, N21,
         N22, N23, N24, N25, N26, N27, n900, n1000, n1100, n120, n130, n140,
         n150, n160, n17, n180, n190, n200, n210, n220, n230, n240, n250, n260,
         n270, n28, n29, n6, n80, n30, n31, n42, n43, n44, n45, n46, n47, n901,
         n91, n92, n93, n94, n96, n99, n1001, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n1101;

  PISO_test_1 PISO_1 ( .out(w2), .in1(in1), .in2(in2), .in3(in3), .in4(in4), 
        .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), 
        .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), 
        .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), 
        .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), 
        .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), 
        .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), 
        .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), 
        .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), 
        .in46(in46), .in47(in47), .in48(in48), .sel(n46), .clk(ex_clk), .rst(
        n44), .test_si(test_si), .test_so(n96), .test_se(n101) );
  counter_PISO_DW01_inc_0 add_107 ( .A(error), .SUM({N27, N26, N25, N24, N23, 
        N22, N21, N20, N19, N18}) );
  counter_PISO_DW01_inc_1 add_104 ( .A(counter), .SUM({N16, N15, N14, N13, N12, 
        N11, N10, N9, N8, N7}) );
  SDFFRQXLTH counter_reg_3_ ( .D(n250), .SI(n109), .SE(n106), .CK(ex_clk), 
        .RN(n44), .Q(counter[3]) );
  SDFFRQXLTH counter_reg_1_ ( .D(n270), .SI(counter[0]), .SE(n107), .CK(ex_clk), .RN(n44), .Q(counter[1]) );
  SDFFRQXLTH counter_reg_2_ ( .D(n260), .SI(n1101), .SE(n105), .CK(ex_clk), 
        .RN(n44), .Q(counter[2]) );
  SDFFRQX1TH counter_reg_9_ ( .D(n200), .SI(counter[8]), .SE(n105), .CK(ex_clk), .RN(n44), .Q(counter[9]) );
  SDFFRQX1TH counter_reg_7_ ( .D(n210), .SI(counter[6]), .SE(n1001), .CK(
        ex_clk), .RN(n44), .Q(counter[7]) );
  SDFFRQX1TH counter_reg_8_ ( .D(n28), .SI(counter[7]), .SE(n1001), .CK(ex_clk), .RN(n44), .Q(counter[8]) );
  SDFFRQX1TH counter_reg_5_ ( .D(n230), .SI(counter[4]), .SE(n99), .CK(ex_clk), 
        .RN(n44), .Q(counter[5]) );
  SDFFRQX1TH counter_reg_4_ ( .D(n240), .SI(n108), .SE(n99), .CK(ex_clk), .RN(
        n44), .Q(counter[4]) );
  SDFFRQX1TH counter_reg_6_ ( .D(n220), .SI(counter[5]), .SE(n106), .CK(ex_clk), .RN(n44), .Q(counter[6]) );
  SDFFRQX1TH counter_reg_0_ ( .D(n29), .SI(n96), .SE(n107), .CK(ex_clk), .RN(
        n44), .Q(counter[0]) );
  SDFFRQX2TH hd_end_reg ( .D(n900), .SI(error[9]), .SE(n105), .CK(ex_clk), 
        .RN(n44), .Q(hd_end) );
  SDFFRQX2TH error_reg_9_ ( .D(n1000), .SI(error[8]), .SE(n105), .CK(ex_clk), 
        .RN(n44), .Q(error[9]) );
  SDFFRQX2TH error_reg_1_ ( .D(n180), .SI(error[0]), .SE(n104), .CK(ex_clk), 
        .RN(n44), .Q(error[1]) );
  SDFFRQX2TH error_reg_2_ ( .D(n17), .SI(error[1]), .SE(n104), .CK(ex_clk), 
        .RN(n44), .Q(error[2]) );
  SDFFRQX2TH error_reg_3_ ( .D(n160), .SI(error[2]), .SE(n107), .CK(ex_clk), 
        .RN(n44), .Q(error[3]) );
  SDFFRQX2TH error_reg_4_ ( .D(n150), .SI(error[3]), .SE(n107), .CK(ex_clk), 
        .RN(n44), .Q(error[4]) );
  SDFFRQX2TH error_reg_5_ ( .D(n140), .SI(error[4]), .SE(n99), .CK(ex_clk), 
        .RN(n44), .Q(error[5]) );
  SDFFRQX2TH error_reg_6_ ( .D(n130), .SI(error[5]), .SE(n106), .CK(ex_clk), 
        .RN(n44), .Q(error[6]) );
  SDFFRQX2TH error_reg_7_ ( .D(n120), .SI(error[6]), .SE(n106), .CK(ex_clk), 
        .RN(n44), .Q(error[7]) );
  SDFFRQX2TH error_reg_8_ ( .D(n1100), .SI(error[7]), .SE(n1001), .CK(ex_clk), 
        .RN(n44), .Q(error[8]) );
  SDFFRQX4TH error_reg_0_ ( .D(n190), .SI(counter[9]), .SE(n103), .CK(ex_clk), 
        .RN(n44), .Q(error[0]) );
  INVX2TH U4 ( .A(1'b1), .Y(out1) );
  CLKAND2X4TH U6 ( .A(n46), .B(n6), .Y(n42) );
  CLKINVX3TH U7 ( .A(n43), .Y(n80) );
  INVX2TH U8 ( .A(n80), .Y(n901) );
  INVXLTH U9 ( .A(counter[0]), .Y(n94) );
  CLKINVX1TH U10 ( .A(n47), .Y(n46) );
  INVXLTH U11 ( .A(w3), .Y(n47) );
  NOR4BX2TH U12 ( .AN(n30), .B(counter[8]), .C(counter[9]), .D(counter[7]), 
        .Y(n6) );
  NAND4XLTH U13 ( .A(n94), .B(n1101), .C(n109), .D(n108), .Y(n31) );
  INVXLTH U14 ( .A(counter[2]), .Y(n93) );
  INVXLTH U15 ( .A(counter[1]), .Y(n92) );
  INVXLTH U16 ( .A(counter[3]), .Y(n91) );
  AO22XLTH U17 ( .A0(error[8]), .A1(n80), .B0(N26), .B1(n901), .Y(n1100) );
  AO22XLTH U18 ( .A0(error[7]), .A1(n80), .B0(N25), .B1(n901), .Y(n120) );
  AO22XLTH U19 ( .A0(error[6]), .A1(n80), .B0(N24), .B1(n901), .Y(n130) );
  AO22XLTH U20 ( .A0(error[5]), .A1(n80), .B0(N23), .B1(n901), .Y(n140) );
  AO22XLTH U21 ( .A0(error[4]), .A1(n80), .B0(N22), .B1(n901), .Y(n150) );
  AO22XLTH U22 ( .A0(error[3]), .A1(n80), .B0(N21), .B1(n901), .Y(n160) );
  AO22XLTH U23 ( .A0(error[2]), .A1(n80), .B0(N20), .B1(n901), .Y(n17) );
  AO22XLTH U24 ( .A0(error[1]), .A1(n80), .B0(N19), .B1(n901), .Y(n180) );
  AO22XLTH U25 ( .A0(error[9]), .A1(n80), .B0(N27), .B1(n901), .Y(n1000) );
  NAND2BXLTH U26 ( .AN(hd_end), .B(n6), .Y(n900) );
  CLKINVX8TH U27 ( .A(n45), .Y(n44) );
  INVXLTH U28 ( .A(rst), .Y(n45) );
  AO22XLTH U29 ( .A0(error[0]), .A1(n80), .B0(N18), .B1(n901), .Y(n190) );
  AO2B2XLTH U30 ( .B0(N11), .B1(n42), .A0(counter[4]), .A1N(n42), .Y(n240) );
  AO2B2XLTH U31 ( .B0(N12), .B1(n42), .A0(counter[5]), .A1N(n42), .Y(n230) );
  OAI2BB2XLTH U32 ( .B0(n42), .B1(n109), .A0N(N9), .A1N(n42), .Y(n260) );
  OAI2BB2XLTH U33 ( .B0(n42), .B1(n1101), .A0N(N8), .A1N(n42), .Y(n270) );
  OAI2BB2XLTH U34 ( .B0(n42), .B1(n108), .A0N(N10), .A1N(n42), .Y(n250) );
  AND2XLTH U36 ( .A(w2), .B(n42), .Y(n43) );
  OAI2BB2XLTH U37 ( .B0(n42), .B1(n94), .A0N(N7), .A1N(n42), .Y(n29) );
  AOI31XLTH U38 ( .A0(counter[4]), .A1(n31), .A2(counter[5]), .B0(counter[6]), 
        .Y(n30) );
  AO21XLTH U39 ( .A0(N13), .A1(n42), .B0(counter[6]), .Y(n220) );
  AO21XLTH U40 ( .A0(N15), .A1(n42), .B0(counter[8]), .Y(n28) );
  AO21XLTH U41 ( .A0(N14), .A1(n42), .B0(counter[7]), .Y(n210) );
  AO21XLTH U42 ( .A0(N16), .A1(n42), .B0(counter[9]), .Y(n200) );
  DLY1X1TH U35 ( .A(test_se), .Y(n99) );
  DLY1X1TH U85 ( .A(test_se), .Y(n1001) );
  DLY1X1TH U86 ( .A(n103), .Y(n101) );
  INVXLTH U87 ( .A(test_se), .Y(n102) );
  INVXLTH U88 ( .A(n102), .Y(n103) );
  INVXLTH U89 ( .A(n102), .Y(n104) );
  DLY1X1TH U90 ( .A(test_se), .Y(n105) );
  DLY1X1TH U91 ( .A(test_se), .Y(n106) );
  DLY1X1TH U92 ( .A(test_se), .Y(n107) );
  DLY1X1TH U93 ( .A(n91), .Y(n108) );
  DLY1X1TH U94 ( .A(n93), .Y(n109) );
  DLY1X1TH U95 ( .A(n92), .Y(n1101) );
endmodule


module fmod2_0 ( out, clk, rst );
  input clk, rst;
  output out;
  wire   n1;

  SDFFRXLTH out_reg ( .D(n1), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst), .Q(out), .QN(n1) );
endmodule


module fmod2_test_0 ( out, clk, rst, test_si, test_se );
  input clk, rst, test_si, test_se;
  output out;
  wire   n1;

  SDFFRXLTH out_reg ( .D(n1), .SI(test_si), .SE(test_se), .CK(clk), .RN(rst), 
        .Q(out), .QN(n1) );
endmodule


module fmod4_test_1 ( out, clk, rst, test_si, test_so, test_se );
  input clk, rst, test_si, test_se;
  output out, test_so;


  fmod2_test_0 f1 ( .out(test_so), .clk(clk), .rst(rst), .test_si(test_si), 
        .test_se(test_se) );
  fmod2_0 f2 ( .out(out), .clk(test_so), .rst(rst) );
endmodule


module sign_xor_23 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25;

  XNOR2X4 U1 ( .A(in1), .B(n5), .Y(n2) );
  CLKXOR2X2 U2 ( .A(in3), .B(in2), .Y(n5) );
  CLKNAND2X12 U3 ( .A(n16), .B(n17), .Y(n1) );
  NAND2X6 U4 ( .A(n2), .B(n3), .Y(n16) );
  CLKNAND2X8 U5 ( .A(n14), .B(n15), .Y(n17) );
  INVX8 U6 ( .A(n2), .Y(n14) );
  INVX6 U7 ( .A(n3), .Y(n15) );
  CLKXOR2X2 U8 ( .A(n4), .B(n23), .Y(n3) );
  XOR2X2 U9 ( .A(in2), .B(n1), .Y(out2) );
  NAND2X2 U11 ( .A(n20), .B(n21), .Y(out1) );
  INVX2 U12 ( .A(n1), .Y(n19) );
  NAND2X1 U13 ( .A(n18), .B(n1), .Y(n21) );
  CLKNAND2X2 U14 ( .A(in1), .B(n19), .Y(n20) );
  XOR2X1 U15 ( .A(n25), .B(n1), .Y(out4) );
  INVXLTH U16 ( .A(in1), .Y(n18) );
  XOR2X1 U17 ( .A(in6), .B(n1), .Y(out6) );
  XOR2XLTH U18 ( .A(in3), .B(n1), .Y(out3) );
  XOR2X3TH U19 ( .A(in6), .B(in5), .Y(n4) );
  XNOR2X1 U10 ( .A(n22), .B(n1), .Y(out5) );
  CLKINVX40 U20 ( .A(in5), .Y(n22) );
  DLY1X1TH U21 ( .A(in4), .Y(n23) );
  INVXLTH U22 ( .A(n23), .Y(n24) );
  INVXLTH U23 ( .A(n24), .Y(n25) );
endmodule


module all6_23 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86;

  sign_xor_23 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  OR2X1 U1 ( .A(n43), .B(n44), .Y(n36) );
  NOR3X4 U3 ( .A(n47), .B(n27), .C(n51), .Y(r6[1]) );
  CLKINVX1 U4 ( .A(n74), .Y(n51) );
  NOR2X4 U5 ( .A(n38), .B(n28), .Y(r5[0]) );
  INVX1TH U6 ( .A(i4[0]), .Y(n50) );
  NOR2X2 U7 ( .A(n36), .B(n28), .Y(r4[0]) );
  OR2X2 U8 ( .A(n54), .B(n63), .Y(n39) );
  NOR3X1 U9 ( .A(n32), .B(n63), .C(n59), .Y(r3[0]) );
  NAND3X2TH U12 ( .A(n71), .B(n69), .C(n67), .Y(n29) );
  NOR2X4 U13 ( .A(n39), .B(n32), .Y(r2[0]) );
  INVX2TH U14 ( .A(i6[0]), .Y(n43) );
  NAND3X3TH U16 ( .A(i5[0]), .B(i4[0]), .C(i6[0]), .Y(n32) );
  OR2XLTH U17 ( .A(n62), .B(n56), .Y(n35) );
  NOR3X1TH U18 ( .A(n65), .B(n57), .C(n52), .Y(r1[2]) );
  OR2X1TH U19 ( .A(n54), .B(n32), .Y(n37) );
  NOR2X2TH U20 ( .A(n35), .B(n29), .Y(r3[3]) );
  INVXLTH U21 ( .A(i1[0]), .Y(n63) );
  CLKINVX1TH U22 ( .A(i2[0]), .Y(n59) );
  NAND3X2TH U23 ( .A(i6[2]), .B(n85), .C(n70), .Y(n30) );
  NOR3X2TH U24 ( .A(n40), .B(n25), .C(n48), .Y(r5[3]) );
  NOR3X2TH U25 ( .A(n41), .B(n26), .C(n78), .Y(r5[2]) );
  NOR3X1TH U26 ( .A(n65), .B(n60), .C(n57), .Y(r3[2]) );
  NOR3X1TH U27 ( .A(n65), .B(n60), .C(n52), .Y(r2[2]) );
  NOR2X3TH U28 ( .A(n37), .B(n59), .Y(r1[0]) );
  OR2X1TH U29 ( .A(n50), .B(n43), .Y(n38) );
  NOR3X4TH U30 ( .A(n31), .B(n61), .C(n58), .Y(r3[1]) );
  INVX2TH U31 ( .A(n73), .Y(n61) );
  NAND3X4TH U32 ( .A(n82), .B(n74), .C(n80), .Y(n31) );
  INVX2TH U33 ( .A(n81), .Y(n58) );
  INVXLTH U34 ( .A(i1[2]), .Y(n60) );
  NOR3X2 U35 ( .A(n31), .B(n58), .C(n79), .Y(r1[1]) );
  NAND3X6 U37 ( .A(i2[0]), .B(i1[0]), .C(i3[0]), .Y(n28) );
  NAND3X4TH U38 ( .A(n81), .B(n73), .C(i3[1]), .Y(n27) );
  NOR3X4TH U39 ( .A(n42), .B(n27), .C(n51), .Y(r5[1]) );
  INVXLTH U40 ( .A(i5[0]), .Y(n44) );
  INVXLTH U41 ( .A(n68), .Y(n62) );
  INVX1TH U42 ( .A(i3[0]), .Y(n54) );
  INVXLTH U43 ( .A(n71), .Y(n45) );
  INVXLTH U45 ( .A(n69), .Y(n48) );
  INVXLTH U46 ( .A(n67), .Y(n40) );
  INVXLTH U47 ( .A(i2[2]), .Y(n57) );
  INVXLTH U48 ( .A(n66), .Y(n55) );
  INVXLTH U49 ( .A(n72), .Y(n56) );
  NOR3X1TH U50 ( .A(n40), .B(n25), .C(n45), .Y(r4[3]) );
  NOR3X1TH U51 ( .A(n45), .B(n25), .C(n48), .Y(r6[3]) );
  NOR3X2 U52 ( .A(n42), .B(n27), .C(n47), .Y(r4[1]) );
  INVXLTH U53 ( .A(n80), .Y(n42) );
  INVX2 U54 ( .A(n82), .Y(n47) );
  NOR3X1TH U55 ( .A(n29), .B(n62), .C(n55), .Y(r2[3]) );
  NOR3X1TH U56 ( .A(n29), .B(n56), .C(n55), .Y(r1[3]) );
  INVXLTH U57 ( .A(i6[2]), .Y(n41) );
  INVXLTH U59 ( .A(n85), .Y(n49) );
  INVXLTH U60 ( .A(i3[2]), .Y(n52) );
  INVXL U61 ( .A(i3[1]), .Y(n53) );
  AND3X8 U2 ( .A(n72), .B(n68), .C(n66), .Y(n64) );
  CLKINVX40 U10 ( .A(n64), .Y(n25) );
  CLKBUFX40 U11 ( .A(n30), .Y(n65) );
  NOR3BX4 U15 ( .AN(i6[2]), .B(n26), .C(n76), .Y(r4[2]) );
  DLY1X1TH U36 ( .A(i3[3]), .Y(n66) );
  DLY1X1TH U44 ( .A(i6[3]), .Y(n67) );
  DLY1X1TH U58 ( .A(i1[3]), .Y(n68) );
  DLY1X1TH U62 ( .A(i4[3]), .Y(n69) );
  DLY1X1TH U63 ( .A(i5[2]), .Y(n70) );
  DLY1X1TH U64 ( .A(i5[3]), .Y(n71) );
  DLY1X1TH U65 ( .A(i2[3]), .Y(n72) );
  DLY1X1TH U66 ( .A(i1[1]), .Y(n73) );
  DLY1X1TH U67 ( .A(i4[1]), .Y(n74) );
  DLY1X1TH U68 ( .A(n70), .Y(n75) );
  INVXLTH U69 ( .A(n75), .Y(n76) );
  INVXLTH U70 ( .A(n75), .Y(n77) );
  INVXLTH U71 ( .A(n85), .Y(n78) );
  INVXLTH U72 ( .A(i3[1]), .Y(n79) );
  DLY1X1TH U73 ( .A(i6[1]), .Y(n80) );
  DLY1X1TH U74 ( .A(i2[1]), .Y(n81) );
  DLY1X1TH U75 ( .A(i5[1]), .Y(n82) );
  NOR3BX4 U76 ( .AN(i5[0]), .B(n28), .C(n50), .Y(r6[0]) );
  AND3X8 U77 ( .A(i2[2]), .B(i1[2]), .C(i3[2]), .Y(n83) );
  CLKINVX40 U78 ( .A(n83), .Y(n26) );
  OR3X8 U79 ( .A(n31), .B(n61), .C(n53), .Y(n84) );
  CLKINVX40 U80 ( .A(n84), .Y(r2[1]) );
  CLKBUFX40 U81 ( .A(i4[2]), .Y(n85) );
  OR3X8 U82 ( .A(n77), .B(n26), .C(n49), .Y(n86) );
  CLKINVX40 U83 ( .A(n86), .Y(r6[2]) );
endmodule


module sign_xor_22 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n14, n15, n16, n17, n18;

  CLKXOR2X2 U1 ( .A(in5), .B(n18), .Y(out5) );
  XOR2X2 U2 ( .A(in3), .B(n18), .Y(out3) );
  XOR2X1 U3 ( .A(in1), .B(n18), .Y(out1) );
  XOR2X3 U4 ( .A(n16), .B(n18), .Y(out6) );
  XOR2X1 U5 ( .A(in2), .B(n18), .Y(out2) );
  XOR2X4 U6 ( .A(n4), .B(in4), .Y(n3) );
  XOR2X2 U7 ( .A(n14), .B(in5), .Y(n4) );
  XNOR2X4TH U8 ( .A(in1), .B(n5), .Y(n2) );
  XOR2X3TH U9 ( .A(in3), .B(in2), .Y(n5) );
  CLKXOR2X2TH U10 ( .A(in4), .B(n18), .Y(out4) );
  XNOR2X4 U11 ( .A(n2), .B(n3), .Y(n1) );
  DLY1X1TH U12 ( .A(in6), .Y(n14) );
  INVXLTH U13 ( .A(n14), .Y(n15) );
  INVXLTH U14 ( .A(n15), .Y(n16) );
  CLKINVX40 U15 ( .A(n1), .Y(n17) );
  CLKINVX40 U16 ( .A(n17), .Y(n18) );
endmodule


module all6_22 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87;

  sign_xor_22 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  INVX1 U1 ( .A(n76), .Y(n66) );
  INVX1 U2 ( .A(n78), .Y(n70) );
  NOR2X2 U3 ( .A(n58), .B(n49), .Y(n41) );
  NOR2X1TH U4 ( .A(n42), .B(n27), .Y(r5[1]) );
  INVX4 U5 ( .A(n41), .Y(n42) );
  INVX2 U6 ( .A(i6[1]), .Y(n49) );
  NAND3X2 U7 ( .A(i3[1]), .B(i1[1]), .C(n75), .Y(n27) );
  INVX2 U8 ( .A(i4[1]), .Y(n58) );
  NOR2X4 U9 ( .A(n43), .B(n28), .Y(r4[0]) );
  INVX2TH U10 ( .A(n87), .Y(n56) );
  NOR3X1 U11 ( .A(n50), .B(n26), .C(n53), .Y(r4[2]) );
  INVX2TH U12 ( .A(n85), .Y(n54) );
  NAND3X4 U13 ( .A(n85), .B(n87), .C(i6[0]), .Y(n32) );
  NOR3X1 U14 ( .A(n53), .B(n26), .C(n59), .Y(r6[2]) );
  NAND3X2 U15 ( .A(i1[2]), .B(n77), .C(n74), .Y(n26) );
  OR2X1TH U16 ( .A(n51), .B(n54), .Y(n43) );
  NAND3X2 U17 ( .A(i3[0]), .B(n78), .C(n76), .Y(n28) );
  INVX2TH U18 ( .A(n46), .Y(n47) );
  NOR2X1TH U19 ( .A(n32), .B(n62), .Y(n46) );
  NOR2X4 U20 ( .A(n47), .B(n66), .Y(r1[0]) );
  INVXLTH U22 ( .A(i6[0]), .Y(n51) );
  NAND3X2TH U23 ( .A(n80), .B(n73), .C(n72), .Y(n25) );
  INVX1TH U24 ( .A(n80), .Y(n67) );
  NAND3X4TH U25 ( .A(n81), .B(n82), .C(i6[3]), .Y(n29) );
  INVX1TH U26 ( .A(n77), .Y(n65) );
  OR2X2TH U27 ( .A(n51), .B(n56), .Y(n44) );
  NOR2X2TH U28 ( .A(n45), .B(n27), .Y(r6[1]) );
  NOR3X4 U29 ( .A(n32), .B(n70), .C(n66), .Y(r3[0]) );
  INVX2TH U30 ( .A(i5[2]), .Y(n53) );
  NOR3X1TH U31 ( .A(n48), .B(n25), .C(n55), .Y(r4[3]) );
  INVXLTH U32 ( .A(n73), .Y(n71) );
  INVXLTH U33 ( .A(i3[1]), .Y(n63) );
  CLKINVX1TH U34 ( .A(n75), .Y(n64) );
  NOR3X4TH U35 ( .A(n30), .B(n68), .C(n65), .Y(r3[2]) );
  OR2XLTH U36 ( .A(n52), .B(n58), .Y(n45) );
  NAND3X3TH U37 ( .A(n79), .B(i4[2]), .C(i5[2]), .Y(n30) );
  INVXLTH U38 ( .A(i3[0]), .Y(n62) );
  NOR3X4TH U39 ( .A(n31), .B(n64), .C(n63), .Y(r1[1]) );
  NAND3X3TH U40 ( .A(i5[1]), .B(i4[1]), .C(i6[1]), .Y(n31) );
  NOR3X4TH U41 ( .A(n49), .B(n27), .C(n52), .Y(r4[1]) );
  NOR2X4TH U42 ( .A(n44), .B(n28), .Y(r5[0]) );
  NOR3X4 U43 ( .A(n30), .B(n65), .C(n61), .Y(r1[2]) );
  INVX2TH U44 ( .A(i5[1]), .Y(n52) );
  NOR3X1TH U45 ( .A(n48), .B(n25), .C(n57), .Y(r5[3]) );
  NOR3X1TH U46 ( .A(n29), .B(n71), .C(n60), .Y(r2[3]) );
  INVXLTH U47 ( .A(n72), .Y(n60) );
  INVXLTH U48 ( .A(i1[2]), .Y(n68) );
  INVXLTH U49 ( .A(i1[1]), .Y(n69) );
  NOR3X4TH U51 ( .A(n31), .B(n69), .C(n64), .Y(r3[1]) );
  NOR3X1 U52 ( .A(n30), .B(n68), .C(n61), .Y(r2[2]) );
  NOR3X2 U53 ( .A(n31), .B(n69), .C(n63), .Y(r2[1]) );
  NOR3X1TH U54 ( .A(n29), .B(n71), .C(n67), .Y(r3[3]) );
  NOR3X1TH U55 ( .A(n29), .B(n67), .C(n60), .Y(r1[3]) );
  NOR3XLTH U56 ( .A(n50), .B(n26), .C(n59), .Y(r5[2]) );
  INVXLTH U57 ( .A(n79), .Y(n50) );
  INVXLTH U58 ( .A(i6[3]), .Y(n48) );
  INVXLTH U59 ( .A(n81), .Y(n55) );
  INVXLTH U60 ( .A(i4[2]), .Y(n59) );
  INVXLTH U61 ( .A(n82), .Y(n57) );
  INVXLTH U62 ( .A(n74), .Y(n61) );
  DLY1X1TH U21 ( .A(i3[3]), .Y(n72) );
  DLY1X1TH U50 ( .A(i1[3]), .Y(n73) );
  DLY1X1TH U63 ( .A(i3[2]), .Y(n74) );
  DLY1X1TH U64 ( .A(i2[1]), .Y(n75) );
  DLY1X1TH U65 ( .A(i2[0]), .Y(n76) );
  DLY1X1TH U66 ( .A(i2[2]), .Y(n77) );
  DLY1X1TH U67 ( .A(i1[0]), .Y(n78) );
  DLY1X1TH U68 ( .A(i6[2]), .Y(n79) );
  DLY1X1TH U69 ( .A(i2[3]), .Y(n80) );
  DLY1X1TH U70 ( .A(i5[3]), .Y(n81) );
  DLY1X1TH U71 ( .A(i4[3]), .Y(n82) );
  INVXLTH U72 ( .A(n55), .Y(n83) );
  OR3X8 U73 ( .A(n54), .B(n28), .C(n56), .Y(n84) );
  CLKINVX40 U74 ( .A(n84), .Y(r6[0]) );
  CLKBUFX40 U75 ( .A(i5[0]), .Y(n85) );
  NOR3BX4 U76 ( .AN(n83), .B(n25), .C(n57), .Y(r6[3]) );
  OR2X8 U77 ( .A(n47), .B(n70), .Y(n86) );
  CLKINVX40 U78 ( .A(n86), .Y(r2[0]) );
  CLKBUFX40 U79 ( .A(i4[0]), .Y(n87) );
endmodule


module sign_xor_21 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n30, n1, n2, n4, n5, n23, n25, n26, n27, n28, n29;

  XOR2XL U1 ( .A(in2), .B(n1), .Y(out2) );
  XOR2X3TH U2 ( .A(in3), .B(in2), .Y(n5) );
  XOR2X1 U3 ( .A(in6), .B(n1), .Y(out6) );
  XOR2X8 U4 ( .A(n2), .B(n23), .Y(n1) );
  XNOR2X4TH U6 ( .A(n26), .B(n5), .Y(n2) );
  XOR2X3TH U7 ( .A(in6), .B(in5), .Y(n4) );
  XOR2XL U8 ( .A(in3), .B(n1), .Y(out3) );
  XOR2X1 U9 ( .A(in5), .B(n1), .Y(n30) );
  XNOR2X4 U10 ( .A(n25), .B(n4), .Y(n23) );
  XOR2X1TH U11 ( .A(n29), .B(n1), .Y(out1) );
  XNOR2X1 U5 ( .A(n27), .B(n1), .Y(out4) );
  CLKBUFX40 U12 ( .A(n30), .Y(out5) );
  DLY1X1TH U13 ( .A(in4), .Y(n25) );
  DLY1X1TH U14 ( .A(in1), .Y(n26) );
  INVXLTH U15 ( .A(n25), .Y(n27) );
  INVXLTH U16 ( .A(n26), .Y(n28) );
  INVXLTH U17 ( .A(n28), .Y(n29) );
endmodule


module all6_21 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86;

  sign_xor_21 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NAND3X2 U1 ( .A(i5[1]), .B(i4[1]), .C(i6[1]), .Y(n31) );
  NOR2X2 U3 ( .A(n53), .B(n57), .Y(n43) );
  NOR2X4 U4 ( .A(n44), .B(n27), .Y(r6[1]) );
  INVX2 U5 ( .A(n43), .Y(n44) );
  NOR2X3 U6 ( .A(n45), .B(n56), .Y(r6[3]) );
  OR2XLTH U7 ( .A(n51), .B(n25), .Y(n45) );
  NOR3X1 U8 ( .A(n49), .B(n26), .C(n52), .Y(r4[2]) );
  NAND3X2 U9 ( .A(i2[0]), .B(i1[0]), .C(i3[0]), .Y(n28) );
  NAND3X2 U10 ( .A(i2[3]), .B(n78), .C(n77), .Y(n25) );
  INVX2 U11 ( .A(n80), .Y(n56) );
  NAND3X2 U12 ( .A(i2[1]), .B(i1[1]), .C(i3[1]), .Y(n27) );
  NOR2X6 U13 ( .A(n46), .B(n58), .Y(r6[0]) );
  NOR3X4 U14 ( .A(n32), .B(n69), .C(n59), .Y(r2[0]) );
  OR2X1TH U16 ( .A(n54), .B(n28), .Y(n46) );
  NOR3X4TH U17 ( .A(n48), .B(n27), .C(n53), .Y(r4[1]) );
  CLKINVX1TH U18 ( .A(i6[1]), .Y(n48) );
  CLKINVX1 U20 ( .A(i1[0]), .Y(n69) );
  NOR3X2 U21 ( .A(n31), .B(n63), .C(n62), .Y(r1[1]) );
  INVXLTH U22 ( .A(i5[0]), .Y(n54) );
  INVXLTH U23 ( .A(i6[2]), .Y(n49) );
  INVX2TH U26 ( .A(i2[0]), .Y(n66) );
  NOR3X1TH U27 ( .A(n30), .B(n70), .C(n65), .Y(r3[2]) );
  INVX1 U28 ( .A(i4[0]), .Y(n58) );
  NOR3X2 U29 ( .A(n50), .B(n28), .C(n54), .Y(r4[0]) );
  INVXLTH U30 ( .A(n74), .Y(n47) );
  INVXLTH U32 ( .A(i6[0]), .Y(n50) );
  INVXLTH U33 ( .A(i3[1]), .Y(n62) );
  NOR3X1TH U34 ( .A(n29), .B(n67), .C(n60), .Y(r2[3]) );
  NOR3X1TH U35 ( .A(n30), .B(n65), .C(n61), .Y(r1[2]) );
  INVX1TH U36 ( .A(i2[1]), .Y(n63) );
  INVXLTH U38 ( .A(n77), .Y(n60) );
  INVXLTH U40 ( .A(n78), .Y(n67) );
  CLKINVX1TH U41 ( .A(i3[0]), .Y(n59) );
  NOR3X1TH U42 ( .A(n29), .B(n64), .C(n60), .Y(r1[3]) );
  NOR3X1TH U43 ( .A(n29), .B(n67), .C(n64), .Y(r3[3]) );
  NOR3X4TH U44 ( .A(n31), .B(n68), .C(n63), .Y(r3[1]) );
  INVXLTH U45 ( .A(i5[3]), .Y(n51) );
  INVXLTH U46 ( .A(i4[2]), .Y(n55) );
  NOR3X1TH U47 ( .A(n47), .B(n25), .C(n51), .Y(r4[3]) );
  INVXLTH U48 ( .A(i2[3]), .Y(n64) );
  NOR3X4TH U50 ( .A(n48), .B(n27), .C(n57), .Y(r5[1]) );
  NOR3X4TH U51 ( .A(n32), .B(n66), .C(n59), .Y(r1[0]) );
  NOR3X2 U53 ( .A(n31), .B(n68), .C(n62), .Y(r2[1]) );
  INVXLTH U54 ( .A(i1[1]), .Y(n68) );
  INVXLTH U55 ( .A(i4[1]), .Y(n57) );
  INVXLTH U56 ( .A(i1[2]), .Y(n70) );
  INVXLTH U57 ( .A(i5[1]), .Y(n53) );
  INVXLTH U58 ( .A(n81), .Y(n52) );
  INVXLTH U59 ( .A(i2[2]), .Y(n65) );
  INVXLTH U60 ( .A(n85), .Y(n61) );
  AND3X8 U2 ( .A(i2[2]), .B(i1[2]), .C(n85), .Y(n71) );
  CLKINVX40 U15 ( .A(n71), .Y(n26) );
  AND3X8 U19 ( .A(i5[3]), .B(n75), .C(n74), .Y(n72) );
  CLKINVX40 U24 ( .A(n72), .Y(n29) );
  NOR3BX4 U25 ( .AN(n74), .B(n25), .C(n56), .Y(r5[3]) );
  NOR3BX4 U31 ( .AN(n82), .B(n70), .C(n61), .Y(r2[2]) );
  OR3X8 U37 ( .A(n32), .B(n69), .C(n66), .Y(n73) );
  CLKINVX40 U39 ( .A(n73), .Y(r3[0]) );
  DLY1X1TH U49 ( .A(i6[3]), .Y(n74) );
  DLY1X1TH U52 ( .A(i4[3]), .Y(n75) );
  INVXLTH U61 ( .A(i4[2]), .Y(n76) );
  DLY1X1TH U62 ( .A(i3[3]), .Y(n77) );
  DLY1X1TH U63 ( .A(i1[3]), .Y(n78) );
  INVXLTH U64 ( .A(n75), .Y(n79) );
  INVXLTH U65 ( .A(n79), .Y(n80) );
  DLY1X1TH U66 ( .A(i5[2]), .Y(n81) );
  NOR3BX4 U67 ( .AN(i6[2]), .B(n26), .C(n76), .Y(r5[2]) );
  NOR3BX4 U68 ( .AN(n81), .B(n26), .C(n55), .Y(r6[2]) );
  AND3X8 U69 ( .A(n81), .B(i4[2]), .C(i6[2]), .Y(n82) );
  CLKINVX40 U70 ( .A(n82), .Y(n30) );
  INVXLTH U71 ( .A(i6[0]), .Y(n83) );
  AND3X8 U72 ( .A(i5[0]), .B(i4[0]), .C(i6[0]), .Y(n84) );
  CLKINVX40 U73 ( .A(n84), .Y(n32) );
  CLKBUFX40 U74 ( .A(i3[2]), .Y(n85) );
  OR3X8 U75 ( .A(n83), .B(n28), .C(n58), .Y(n86) );
  CLKINVX40 U76 ( .A(n86), .Y(r5[0]) );
endmodule


module sign_xor_20 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n4, n5, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50;

  NAND2X2 U1 ( .A(n41), .B(n42), .Y(out1) );
  CLKINVX24 U2 ( .A(n1), .Y(n37) );
  BUFX8 U3 ( .A(in4), .Y(n35) );
  CLKNAND2X2 U4 ( .A(n44), .B(n45), .Y(out5) );
  NAND2XL U5 ( .A(in1), .B(n37), .Y(n41) );
  NAND2XLTH U6 ( .A(n35), .B(n37), .Y(n38) );
  NAND2XLTH U7 ( .A(n36), .B(n1), .Y(n39) );
  CLKNAND2X4 U8 ( .A(n38), .B(n39), .Y(out4) );
  INVXLTH U9 ( .A(n35), .Y(n36) );
  XOR2XL U10 ( .A(in3), .B(n1), .Y(out3) );
  NAND2XLTH U11 ( .A(n40), .B(n1), .Y(n42) );
  XOR2X1TH U12 ( .A(in6), .B(n1), .Y(out6) );
  XOR2X1TH U13 ( .A(in2), .B(n1), .Y(out2) );
  INVX6 U14 ( .A(n2), .Y(n46) );
  INVXLTH U15 ( .A(in1), .Y(n40) );
  NAND2X3 U16 ( .A(n46), .B(n50), .Y(n49) );
  XOR2X2TH U17 ( .A(in6), .B(in5), .Y(n4) );
  XOR2X3TH U18 ( .A(in3), .B(in2), .Y(n5) );
  NAND2XLTH U19 ( .A(in5), .B(n37), .Y(n44) );
  NAND2XLTH U20 ( .A(n43), .B(n1), .Y(n45) );
  INVXLTH U21 ( .A(in5), .Y(n43) );
  NAND2X4 U22 ( .A(n2), .B(n47), .Y(n48) );
  INVX4 U23 ( .A(n50), .Y(n47) );
  NAND2X8 U24 ( .A(n48), .B(n49), .Y(n1) );
  XNOR2X4 U25 ( .A(in1), .B(n5), .Y(n2) );
  XNOR2X4 U26 ( .A(n35), .B(n4), .Y(n50) );
endmodule


module all6_20 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93;

  sign_xor_20 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR2X2 U1 ( .A(n52), .B(n28), .Y(r5[0]) );
  NOR3X1 U2 ( .A(n30), .B(n77), .C(n69), .Y(r2[2]) );
  NAND3X4 U3 ( .A(n85), .B(i4[2]), .C(i5[2]), .Y(n30) );
  NAND3X2 U5 ( .A(n84), .B(n81), .C(n82), .Y(n29) );
  NOR2X1 U6 ( .A(n64), .B(n62), .Y(n50) );
  NOR2X4 U7 ( .A(n51), .B(n28), .Y(r6[0]) );
  INVX2 U8 ( .A(n50), .Y(n51) );
  INVXLTH U9 ( .A(i5[0]), .Y(n62) );
  NAND2X6 U10 ( .A(i3[0]), .B(n53), .Y(n28) );
  INVXLTH U11 ( .A(i4[0]), .Y(n64) );
  NOR2X4TH U13 ( .A(n54), .B(n74), .Y(r3[0]) );
  OR2X2TH U14 ( .A(n57), .B(n64), .Y(n52) );
  NOR3X4 U15 ( .A(n32), .B(n75), .C(n70), .Y(r2[0]) );
  NAND3X4 U16 ( .A(i5[0]), .B(i4[0]), .C(i6[0]), .Y(n32) );
  NOR3X4 U17 ( .A(n58), .B(n27), .C(n61), .Y(r4[1]) );
  NOR3X4 U18 ( .A(n57), .B(n28), .C(n62), .Y(r4[0]) );
  NOR3X2TH U19 ( .A(n29), .B(n78), .C(n73), .Y(r3[3]) );
  INVX2TH U21 ( .A(i3[0]), .Y(n70) );
  CLKINVX1TH U22 ( .A(i2[0]), .Y(n74) );
  NOR3X1TH U23 ( .A(n60), .B(n26), .C(n87), .Y(r6[2]) );
  INVX2TH U24 ( .A(i6[1]), .Y(n58) );
  INVX1TH U25 ( .A(n83), .Y(n76) );
  INVX1TH U26 ( .A(i3[1]), .Y(n67) );
  NAND3X4TH U27 ( .A(i5[1]), .B(i4[1]), .C(i6[1]), .Y(n31) );
  NOR3X1TH U28 ( .A(n30), .B(n72), .C(n69), .Y(r1[2]) );
  NOR3X1TH U29 ( .A(n30), .B(n77), .C(n72), .Y(r3[2]) );
  INVX2 U30 ( .A(i4[1]), .Y(n66) );
  NAND3X2 U31 ( .A(i2[3]), .B(i1[3]), .C(i3[3]), .Y(n25) );
  NOR3X4 U32 ( .A(n32), .B(n74), .C(n70), .Y(r1[0]) );
  NOR3X4 U33 ( .A(n31), .B(n71), .C(n67), .Y(r1[1]) );
  NOR3X4 U34 ( .A(n56), .B(n26), .C(n60), .Y(r4[2]) );
  NOR3X4TH U35 ( .A(n31), .B(n76), .C(n71), .Y(r3[1]) );
  INVX2TH U36 ( .A(i1[0]), .Y(n75) );
  INVXLTH U37 ( .A(i2[2]), .Y(n72) );
  CLKINVX1TH U38 ( .A(i2[1]), .Y(n71) );
  AND2XLTH U40 ( .A(i1[0]), .B(i2[0]), .Y(n53) );
  OR2XLTH U41 ( .A(n75), .B(n32), .Y(n54) );
  NOR3X4TH U42 ( .A(n55), .B(n25), .C(n89), .Y(r4[3]) );
  NAND3X2TH U43 ( .A(i2[2]), .B(i1[2]), .C(i3[2]), .Y(n26) );
  INVXLTH U44 ( .A(i1[3]), .Y(n78) );
  INVXLTH U45 ( .A(i1[2]), .Y(n77) );
  INVXLTH U46 ( .A(i2[3]), .Y(n73) );
  NOR3X1TH U48 ( .A(n55), .B(n25), .C(n65), .Y(r5[3]) );
  CLKINVX1TH U50 ( .A(i6[0]), .Y(n57) );
  INVXLTH U51 ( .A(i3[2]), .Y(n69) );
  INVXLTH U54 ( .A(i5[1]), .Y(n61) );
  INVXLTH U55 ( .A(n85), .Y(n56) );
  INVXLTH U56 ( .A(n82), .Y(n55) );
  INVXLTH U57 ( .A(i5[2]), .Y(n60) );
  INVXLTH U58 ( .A(n84), .Y(n59) );
  INVXLTH U59 ( .A(i4[2]), .Y(n63) );
  INVXLTH U60 ( .A(n81), .Y(n65) );
  AND3X8 U4 ( .A(i2[1]), .B(n83), .C(i3[1]), .Y(n79) );
  CLKINVX40 U12 ( .A(n79), .Y(n27) );
  NOR3BX4 U20 ( .AN(i6[1]), .B(n27), .C(n66), .Y(r5[1]) );
  NOR3BX4 U39 ( .AN(i5[1]), .B(n27), .C(n66), .Y(r6[1]) );
  NAND3BX4 U47 ( .AN(n29), .B(i2[3]), .C(i3[3]), .Y(n80) );
  CLKINVX40 U49 ( .A(n80), .Y(r1[3]) );
  DLY1X1TH U52 ( .A(i4[3]), .Y(n81) );
  DLY1X1TH U53 ( .A(i6[3]), .Y(n82) );
  DLY1X1TH U61 ( .A(i1[1]), .Y(n83) );
  DLY1X1TH U62 ( .A(i5[3]), .Y(n84) );
  DLY1X1TH U63 ( .A(i6[2]), .Y(n85) );
  DLY1X1TH U64 ( .A(n65), .Y(n86) );
  INVXLTH U65 ( .A(i4[2]), .Y(n87) );
  DLY1X1TH U66 ( .A(n56), .Y(n88) );
  DLY1X1TH U67 ( .A(n59), .Y(n89) );
  NAND3BX4 U68 ( .AN(n29), .B(i1[3]), .C(i3[3]), .Y(n90) );
  CLKINVX40 U69 ( .A(n90), .Y(r2[3]) );
  OR3X8 U70 ( .A(n76), .B(n31), .C(n67), .Y(n91) );
  CLKINVX40 U71 ( .A(n91), .Y(r2[1]) );
  OR3X8 U72 ( .A(n88), .B(n26), .C(n63), .Y(n92) );
  CLKINVX40 U73 ( .A(n92), .Y(r5[2]) );
  OR3X8 U74 ( .A(n89), .B(n25), .C(n86), .Y(n93) );
  CLKINVX40 U75 ( .A(n93), .Y(r6[3]) );
endmodule


module sign_xor_19 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25;

  XOR2XLTH U1 ( .A(n23), .B(n1), .Y(out1) );
  XOR2X3 U2 ( .A(in3), .B(in2), .Y(n5) );
  CLKXOR2X4 U3 ( .A(n4), .B(n21), .Y(n3) );
  XOR2X3 U4 ( .A(in6), .B(in5), .Y(n4) );
  CLKNAND2X4 U5 ( .A(in3), .B(n12), .Y(n13) );
  NAND2XLTH U6 ( .A(n11), .B(n1), .Y(n14) );
  NAND2X4 U7 ( .A(n13), .B(n14), .Y(out3) );
  INVXLTH U8 ( .A(in3), .Y(n11) );
  INVXLTH U9 ( .A(n1), .Y(n12) );
  CLKNAND2X12 U10 ( .A(n17), .B(n18), .Y(n1) );
  NAND2X4 U11 ( .A(n2), .B(n3), .Y(n17) );
  NAND2X5 U12 ( .A(n15), .B(n16), .Y(n18) );
  INVX6 U13 ( .A(n2), .Y(n15) );
  CLKINVX4 U14 ( .A(n3), .Y(n16) );
  XNOR2X2 U15 ( .A(n20), .B(n5), .Y(n2) );
  XOR2XLTH U17 ( .A(in5), .B(n1), .Y(out5) );
  XOR2XLTH U18 ( .A(n25), .B(n1), .Y(out4) );
  XOR2X1 U19 ( .A(in6), .B(n1), .Y(out6) );
  XNOR2X1 U16 ( .A(n19), .B(n1), .Y(out2) );
  CLKINVX40 U20 ( .A(in2), .Y(n19) );
  DLY1X1TH U21 ( .A(in1), .Y(n20) );
  DLY1X1TH U22 ( .A(in4), .Y(n21) );
  INVXLTH U23 ( .A(n20), .Y(n22) );
  INVXLTH U24 ( .A(n22), .Y(n23) );
  INVXLTH U25 ( .A(n21), .Y(n24) );
  INVXLTH U26 ( .A(n24), .Y(n25) );
endmodule


module all6_19 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n41, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82;

  NOR3X1 U50 ( .A(n30), .B(n67), .C(n59), .Y(r2[2]) );
  sign_xor_19 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  INVX2 U1 ( .A(i1[0]), .Y(n66) );
  NOR3X1 U2 ( .A(n29), .B(n69), .C(n61), .Y(r2[3]) );
  NOR2X2 U3 ( .A(n52), .B(n57), .Y(n41) );
  NOR2X4 U7 ( .A(n45), .B(n32), .Y(r2[0]) );
  NOR2X2TH U8 ( .A(n43), .B(n25), .Y(r6[3]) );
  NAND3X2 U9 ( .A(i5[1]), .B(n76), .C(n72), .Y(n31) );
  NOR3X4TH U10 ( .A(n32), .B(n65), .C(n58), .Y(r1[0]) );
  NOR3X1 U11 ( .A(n47), .B(n26), .C(n55), .Y(r5[2]) );
  OR2XLTH U12 ( .A(n54), .B(n53), .Y(n43) );
  NOR3X1 U13 ( .A(n29), .B(n69), .C(n64), .Y(r3[3]) );
  NOR3X2 U14 ( .A(n48), .B(n27), .C(n56), .Y(r5[1]) );
  NAND3X2 U15 ( .A(n74), .B(n73), .C(n71), .Y(n25) );
  NOR3X1 U16 ( .A(n30), .B(n62), .C(n59), .Y(r1[2]) );
  NOR3X1TH U17 ( .A(n49), .B(n25), .C(n54), .Y(r5[3]) );
  NOR3X1TH U18 ( .A(n30), .B(n67), .C(n62), .Y(r3[2]) );
  OR2X1TH U19 ( .A(n66), .B(n58), .Y(n45) );
  INVXL U20 ( .A(i2[1]), .Y(n63) );
  OR2X1 U21 ( .A(n70), .B(n63), .Y(n44) );
  NAND3X2TH U22 ( .A(i5[3]), .B(i4[3]), .C(n78), .Y(n29) );
  INVX1TH U23 ( .A(i3[0]), .Y(n58) );
  INVX1TH U24 ( .A(n82), .Y(n68) );
  INVXLTH U25 ( .A(n77), .Y(n60) );
  NOR3X4TH U26 ( .A(n29), .B(n64), .C(n61), .Y(r1[3]) );
  NAND3X3 U27 ( .A(n75), .B(i1[2]), .C(i3[2]), .Y(n26) );
  CLKINVX1 U28 ( .A(i2[0]), .Y(n65) );
  NOR2X4 U29 ( .A(n44), .B(n31), .Y(r1[1]) );
  NOR3X1 U30 ( .A(n46), .B(n28), .C(n57), .Y(r5[0]) );
  INVX1TH U31 ( .A(i4[0]), .Y(n57) );
  NAND3X4TH U32 ( .A(n77), .B(n82), .C(i2[1]), .Y(n27) );
  INVXLTH U33 ( .A(i5[1]), .Y(n51) );
  NOR3X1TH U34 ( .A(n50), .B(n26), .C(n55), .Y(r6[2]) );
  INVX1TH U35 ( .A(i5[0]), .Y(n52) );
  INVXLTH U37 ( .A(n71), .Y(n61) );
  INVXLTH U38 ( .A(n74), .Y(n64) );
  NAND3X4TH U39 ( .A(i5[0]), .B(i4[0]), .C(i6[0]), .Y(n32) );
  INVX2TH U40 ( .A(n76), .Y(n56) );
  INVXLTH U41 ( .A(n78), .Y(n49) );
  INVXLTH U42 ( .A(i4[3]), .Y(n54) );
  INVXLTH U43 ( .A(i5[3]), .Y(n53) );
  INVXLTH U45 ( .A(n73), .Y(n69) );
  INVXLTH U46 ( .A(n72), .Y(n48) );
  NOR3X1TH U47 ( .A(n49), .B(n25), .C(n53), .Y(r4[3]) );
  NAND3X2TH U48 ( .A(i5[2]), .B(i4[2]), .C(i6[2]), .Y(n30) );
  INVXLTH U49 ( .A(i6[0]), .Y(n46) );
  NOR3X4 U52 ( .A(n32), .B(n66), .C(n65), .Y(r3[0]) );
  NOR3X4TH U54 ( .A(n31), .B(n68), .C(n63), .Y(r3[1]) );
  NOR3XLTH U55 ( .A(n47), .B(n26), .C(n50), .Y(r4[2]) );
  INVXLTH U56 ( .A(i6[2]), .Y(n47) );
  INVXLTH U57 ( .A(i1[2]), .Y(n67) );
  INVXLTH U58 ( .A(i5[2]), .Y(n50) );
  INVXLTH U59 ( .A(n75), .Y(n62) );
  INVXLTH U60 ( .A(i4[2]), .Y(n55) );
  INVXLTH U61 ( .A(i3[2]), .Y(n59) );
  NOR3BX4 U4 ( .AN(i5[1]), .B(n27), .C(n56), .Y(r6[1]) );
  INVXLTH U5 ( .A(n77), .Y(n70) );
  DLY1X1TH U6 ( .A(i3[3]), .Y(n71) );
  DLY1X1TH U36 ( .A(i6[1]), .Y(n72) );
  DLY1X1TH U44 ( .A(i1[3]), .Y(n73) );
  DLY1X1TH U51 ( .A(i2[3]), .Y(n74) );
  DLY1X1TH U53 ( .A(i2[2]), .Y(n75) );
  DLY1X1TH U62 ( .A(i4[1]), .Y(n76) );
  DLY1X1TH U63 ( .A(i3[1]), .Y(n77) );
  DLY1X1TH U64 ( .A(i6[3]), .Y(n78) );
  INVXLTH U65 ( .A(n48), .Y(n79) );
  OR3X8 U66 ( .A(n60), .B(n68), .C(n31), .Y(n80) );
  CLKINVX40 U67 ( .A(n80), .Y(r2[1]) );
  AND2X8 U68 ( .A(n41), .B(n81), .Y(r6[0]) );
  AND3X8 U69 ( .A(i2[0]), .B(i1[0]), .C(i3[0]), .Y(n81) );
  CLKINVX40 U70 ( .A(n81), .Y(n28) );
  NOR3BX4 U71 ( .AN(i6[0]), .B(n28), .C(n52), .Y(r4[0]) );
  CLKBUFX40 U72 ( .A(i1[1]), .Y(n82) );
  NOR3BX4 U73 ( .AN(n79), .B(n27), .C(n51), .Y(r4[1]) );
endmodule


module sign_xor_18 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n4, n5, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25;

  XOR2X8 U1 ( .A(n2), .B(n18), .Y(n1) );
  XOR2X2 U2 ( .A(in3), .B(in2), .Y(n5) );
  INVX2TH U3 ( .A(n25), .Y(n15) );
  CLKNAND2X2 U4 ( .A(in1), .B(n15), .Y(n12) );
  NAND2XLTH U5 ( .A(n11), .B(n25), .Y(n13) );
  NAND2X2 U6 ( .A(n12), .B(n13), .Y(out1) );
  INVXLTH U7 ( .A(in1), .Y(n11) );
  XOR2X1 U9 ( .A(in5), .B(n25), .Y(out5) );
  NAND2X1 U10 ( .A(in2), .B(n15), .Y(n16) );
  XOR2X1 U12 ( .A(in3), .B(n25), .Y(out3) );
  INVXLTH U13 ( .A(in2), .Y(n14) );
  XOR2X4TH U15 ( .A(in6), .B(in5), .Y(n4) );
  XNOR2X4TH U16 ( .A(in1), .B(n5), .Y(n2) );
  XOR2X1TH U17 ( .A(n23), .B(n25), .Y(out4) );
  XNOR2X4 U18 ( .A(n21), .B(n4), .Y(n18) );
  XNOR2X1 U8 ( .A(in6), .B(n24), .Y(out6) );
  AND2X8 U11 ( .A(n14), .B(n25), .Y(n19) );
  CLKINVX40 U14 ( .A(n19), .Y(n17) );
  AND2X8 U19 ( .A(n16), .B(n17), .Y(n20) );
  CLKINVX40 U20 ( .A(n20), .Y(out2) );
  DLY1X1TH U21 ( .A(in4), .Y(n21) );
  INVXLTH U22 ( .A(n21), .Y(n22) );
  INVXLTH U23 ( .A(n22), .Y(n23) );
  CLKINVX40 U24 ( .A(n1), .Y(n24) );
  CLKINVX40 U25 ( .A(n24), .Y(n25) );
endmodule


module all6_18 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86;

  NOR3X1 U34 ( .A(n57), .B(n26), .C(n60), .Y(r6[2]) );
  sign_xor_18 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NAND3X3 U1 ( .A(i5[0]), .B(i4[0]), .C(i6[0]), .Y(n32) );
  NAND3X3 U2 ( .A(n84), .B(i2[0]), .C(i3[0]), .Y(n28) );
  NOR2X4 U3 ( .A(n46), .B(n32), .Y(r1[0]) );
  NOR2X4TH U4 ( .A(n49), .B(n28), .Y(r6[0]) );
  NOR3X4 U5 ( .A(n56), .B(n27), .C(n61), .Y(r6[1]) );
  NOR3X4TH U6 ( .A(n51), .B(n27), .C(n56), .Y(r4[1]) );
  NOR3X2 U7 ( .A(n51), .B(n27), .C(n61), .Y(r5[1]) );
  NAND2X2 U8 ( .A(i1[1]), .B(n47), .Y(n27) );
  NOR3X4 U9 ( .A(n52), .B(n28), .C(n59), .Y(r5[0]) );
  NOR3X1 U10 ( .A(n52), .B(n28), .C(n55), .Y(r4[0]) );
  INVX2 U11 ( .A(i5[0]), .Y(n55) );
  NOR3X2 U12 ( .A(n30), .B(n69), .C(n62), .Y(r1[2]) );
  NAND3X4 U13 ( .A(i5[1]), .B(i4[1]), .C(i6[1]), .Y(n31) );
  NAND3X4 U14 ( .A(i5[2]), .B(i4[2]), .C(i6[2]), .Y(n30) );
  OR2XLTH U15 ( .A(n30), .B(n62), .Y(n45) );
  OR2XLTH U16 ( .A(n64), .B(n67), .Y(n46) );
  INVX2TH U17 ( .A(i4[0]), .Y(n59) );
  INVX2TH U18 ( .A(n84), .Y(n70) );
  NOR3X1TH U19 ( .A(n53), .B(n25), .C(n58), .Y(r5[3]) );
  INVX1TH U20 ( .A(i1[1]), .Y(n71) );
  AND2XLTH U21 ( .A(i3[1]), .B(i2[1]), .Y(n47) );
  NAND3X3 U22 ( .A(n81), .B(i2[2]), .C(i3[2]), .Y(n26) );
  OR2X2TH U23 ( .A(n55), .B(n59), .Y(n49) );
  NOR2X4 U24 ( .A(n45), .B(n73), .Y(r2[2]) );
  INVX2 U25 ( .A(i3[2]), .Y(n62) );
  INVXLTH U26 ( .A(n81), .Y(n73) );
  INVX1TH U27 ( .A(i3[0]), .Y(n64) );
  CLKINVX1TH U28 ( .A(i4[1]), .Y(n61) );
  CLKINVX1TH U29 ( .A(i5[1]), .Y(n56) );
  CLKINVX1TH U30 ( .A(i6[0]), .Y(n52) );
  INVXLTH U31 ( .A(i2[2]), .Y(n69) );
  NOR3X2TH U32 ( .A(n29), .B(n72), .C(n63), .Y(r2[3]) );
  NOR2X2TH U33 ( .A(n48), .B(n65), .Y(r2[1]) );
  OR2XLTH U35 ( .A(n31), .B(n71), .Y(n48) );
  NOR3X1TH U36 ( .A(n31), .B(n71), .C(n68), .Y(r3[1]) );
  NOR3X1TH U37 ( .A(n30), .B(n73), .C(n69), .Y(r3[2]) );
  INVXLTH U38 ( .A(n76), .Y(n53) );
  NAND3X2TH U39 ( .A(n80), .B(n77), .C(n75), .Y(n25) );
  INVXLTH U40 ( .A(n79), .Y(n54) );
  NOR3X1TH U41 ( .A(n53), .B(n25), .C(n54), .Y(r4[3]) );
  NOR3X1TH U42 ( .A(n54), .B(n25), .C(n58), .Y(r6[3]) );
  NOR3X1TH U43 ( .A(n29), .B(n66), .C(n63), .Y(r1[3]) );
  NOR3X4TH U44 ( .A(n31), .B(n68), .C(n65), .Y(r1[1]) );
  INVXLTH U45 ( .A(n78), .Y(n58) );
  INVXLTH U46 ( .A(i2[0]), .Y(n67) );
  INVXLTH U47 ( .A(i4[2]), .Y(n60) );
  INVXLTH U48 ( .A(i6[2]), .Y(n50) );
  INVXLTH U49 ( .A(i5[2]), .Y(n57) );
  CLKINVX1TH U50 ( .A(i6[1]), .Y(n51) );
  INVXLTH U51 ( .A(n77), .Y(n72) );
  INVXLTH U53 ( .A(n80), .Y(n66) );
  INVXLTH U54 ( .A(n75), .Y(n63) );
  NOR3X1TH U55 ( .A(n29), .B(n72), .C(n66), .Y(r3[3]) );
  NOR3XLTH U56 ( .A(n50), .B(n26), .C(n57), .Y(r4[2]) );
  NOR3X4TH U58 ( .A(n32), .B(n70), .C(n67), .Y(r3[0]) );
  INVXLTH U60 ( .A(i2[1]), .Y(n68) );
  INVXLTH U61 ( .A(i3[1]), .Y(n65) );
  AND3X8 U52 ( .A(n79), .B(n78), .C(n76), .Y(n74) );
  CLKINVX40 U57 ( .A(n74), .Y(n29) );
  DLY1X1TH U59 ( .A(i3[3]), .Y(n75) );
  DLY1X1TH U62 ( .A(i6[3]), .Y(n76) );
  DLY1X1TH U63 ( .A(i1[3]), .Y(n77) );
  DLY1X1TH U64 ( .A(i4[3]), .Y(n78) );
  DLY1X1TH U65 ( .A(i5[3]), .Y(n79) );
  DLY1X1TH U66 ( .A(i2[3]), .Y(n80) );
  DLY1X1TH U67 ( .A(i1[2]), .Y(n81) );
  DLY1X1TH U68 ( .A(n50), .Y(n82) );
  DLY1X1TH U69 ( .A(n60), .Y(n83) );
  DLY1X1TH U70 ( .A(i1[0]), .Y(n84) );
  OR3X8 U71 ( .A(n32), .B(n70), .C(n64), .Y(n85) );
  CLKINVX40 U72 ( .A(n85), .Y(r2[0]) );
  OR3X8 U73 ( .A(n82), .B(n26), .C(n83), .Y(n86) );
  CLKINVX40 U74 ( .A(n86), .Y(r5[2]) );
endmodule


module sign_xor_17 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n4, n5, n26, n27, n28, n29, n30, n31, n32, n33;

  INVXLTH U1 ( .A(n1), .Y(n27) );
  NAND2X2 U2 ( .A(n28), .B(n29), .Y(out4) );
  XOR2XLTH U3 ( .A(in6), .B(n1), .Y(out6) );
  NAND2XLTH U4 ( .A(in4), .B(n27), .Y(n28) );
  NAND2XLTH U5 ( .A(n26), .B(n1), .Y(n29) );
  INVXLTH U6 ( .A(in4), .Y(n26) );
  CLKXOR2X12 U7 ( .A(n2), .B(n30), .Y(n1) );
  XOR2XLTH U8 ( .A(in3), .B(n1), .Y(out3) );
  XOR2X4TH U9 ( .A(in3), .B(in2), .Y(n5) );
  XOR2X2TH U10 ( .A(in6), .B(in5), .Y(n4) );
  XOR2X1TH U11 ( .A(n33), .B(n1), .Y(out1) );
  XNOR2X4TH U12 ( .A(n31), .B(n5), .Y(n2) );
  XOR2X1TH U13 ( .A(in2), .B(n1), .Y(out2) );
  XNOR2X4 U14 ( .A(in4), .B(n4), .Y(n30) );
  XOR2X1TH U15 ( .A(in5), .B(n1), .Y(out5) );
  DLY1X1TH U16 ( .A(in1), .Y(n31) );
  INVXLTH U17 ( .A(n31), .Y(n32) );
  INVXLTH U18 ( .A(n32), .Y(n33) );
endmodule


module all6_17 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85;

  NAND3X2 U2 ( .A(i3[2]), .B(i1[2]), .C(n76), .Y(n26) );
  sign_xor_17 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X1 U1 ( .A(n29), .B(n67), .C(n64), .Y(r1[3]) );
  INVXL U3 ( .A(n76), .Y(n65) );
  AND2XLTH U5 ( .A(i6[0]), .B(i5[0]), .Y(n48) );
  NOR3X4 U6 ( .A(n32), .B(n72), .C(n63), .Y(r2[0]) );
  NAND3X4 U7 ( .A(n77), .B(i1[1]), .C(n84), .Y(n27) );
  INVXL U8 ( .A(i6[1]), .Y(n52) );
  NAND2X2 U9 ( .A(i4[0]), .B(n48), .Y(n32) );
  CLKINVX1 U10 ( .A(i4[0]), .Y(n60) );
  NOR3X4 U11 ( .A(n56), .B(n28), .C(n60), .Y(r6[0]) );
  INVX1 U12 ( .A(i5[0]), .Y(n56) );
  CLKINVX1 U13 ( .A(n81), .Y(n63) );
  CLKINVX1 U14 ( .A(n78), .Y(n68) );
  NOR3X1TH U15 ( .A(n29), .B(n70), .C(n64), .Y(r2[3]) );
  CLKINVX1TH U16 ( .A(n80), .Y(n72) );
  INVXLTH U17 ( .A(n84), .Y(n62) );
  NAND3X2TH U18 ( .A(i5[1]), .B(i4[1]), .C(i6[1]), .Y(n31) );
  NOR3X2TH U19 ( .A(n50), .B(n26), .C(n53), .Y(r4[2]) );
  NOR3X1TH U20 ( .A(n30), .B(n69), .C(n65), .Y(r3[2]) );
  NOR3X4 U21 ( .A(n31), .B(n66), .C(n62), .Y(r1[1]) );
  NOR3X4 U22 ( .A(n32), .B(n72), .C(n68), .Y(r3[0]) );
  NOR3X2 U23 ( .A(n31), .B(n71), .C(n62), .Y(r2[1]) );
  NAND3X2TH U24 ( .A(i2[3]), .B(i1[3]), .C(i3[3]), .Y(n25) );
  INVXLTH U25 ( .A(n75), .Y(n49) );
  INVXLTH U26 ( .A(i1[3]), .Y(n70) );
  NAND3X2TH U27 ( .A(i5[3]), .B(i4[3]), .C(n75), .Y(n29) );
  INVXLTH U28 ( .A(i2[3]), .Y(n67) );
  INVXLTH U29 ( .A(n77), .Y(n66) );
  NOR3X1TH U30 ( .A(n53), .B(n26), .C(n58), .Y(r6[2]) );
  INVXLTH U31 ( .A(i4[2]), .Y(n58) );
  NAND3X4 U32 ( .A(n79), .B(i4[2]), .C(i6[2]), .Y(n30) );
  NOR3X4TH U33 ( .A(n54), .B(n27), .C(n82), .Y(r6[1]) );
  NOR3X4 U34 ( .A(n30), .B(n65), .C(n61), .Y(r1[2]) );
  INVXLTH U36 ( .A(i5[3]), .Y(n55) );
  INVXLTH U37 ( .A(i3[3]), .Y(n64) );
  NOR3X1TH U38 ( .A(n55), .B(n25), .C(n57), .Y(r6[3]) );
  NOR3X1TH U39 ( .A(n49), .B(n25), .C(n55), .Y(r4[3]) );
  INVXLTH U40 ( .A(i4[3]), .Y(n57) );
  NOR3X1TH U41 ( .A(n49), .B(n25), .C(n57), .Y(r5[3]) );
  INVXLTH U42 ( .A(n79), .Y(n53) );
  NOR3X1TH U43 ( .A(n29), .B(n70), .C(n67), .Y(r3[3]) );
  INVXLTH U44 ( .A(i1[1]), .Y(n71) );
  NOR3X2TH U45 ( .A(n31), .B(n71), .C(n66), .Y(r3[1]) );
  CLKINVX1TH U46 ( .A(i6[0]), .Y(n51) );
  NOR3X2 U47 ( .A(n74), .B(n27), .C(n54), .Y(r4[1]) );
  NOR3XLTH U49 ( .A(n30), .B(n69), .C(n61), .Y(r2[2]) );
  NAND3X4 U50 ( .A(n78), .B(n80), .C(n81), .Y(n28) );
  INVX2 U51 ( .A(i6[2]), .Y(n50) );
  INVXLTH U52 ( .A(i1[2]), .Y(n69) );
  INVXLTH U53 ( .A(i5[1]), .Y(n54) );
  INVXLTH U54 ( .A(i4[1]), .Y(n59) );
  INVXLTH U55 ( .A(i3[2]), .Y(n61) );
  NOR3X4TH U56 ( .A(n51), .B(n28), .C(n56), .Y(r4[0]) );
  NOR3X4TH U57 ( .A(n51), .B(n28), .C(n60), .Y(r5[0]) );
  OR3X8 U4 ( .A(n32), .B(n68), .C(n63), .Y(n73) );
  CLKINVX40 U35 ( .A(n73), .Y(r1[0]) );
  INVXLTH U48 ( .A(i6[1]), .Y(n74) );
  DLY1X1TH U58 ( .A(i6[3]), .Y(n75) );
  DLY1X1TH U59 ( .A(i2[2]), .Y(n76) );
  DLY1X1TH U60 ( .A(i2[1]), .Y(n77) );
  DLY1X1TH U61 ( .A(i2[0]), .Y(n78) );
  DLY1X1TH U62 ( .A(i5[2]), .Y(n79) );
  DLY1X1TH U63 ( .A(i1[0]), .Y(n80) );
  DLY1X1TH U64 ( .A(i3[0]), .Y(n81) );
  INVXLTH U65 ( .A(i4[1]), .Y(n82) );
  OR3X8 U66 ( .A(n52), .B(n27), .C(n59), .Y(n83) );
  CLKINVX40 U67 ( .A(n83), .Y(r5[1]) );
  CLKBUFX40 U68 ( .A(i3[1]), .Y(n84) );
  NOR3BX4 U69 ( .AN(n85), .B(n26), .C(n58), .Y(r5[2]) );
  CLKINVX40 U70 ( .A(n50), .Y(n85) );
endmodule


module sign_xor_16 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48;

  NAND2X2TH U1 ( .A(in6), .B(n32), .Y(n33) );
  NAND2XLTH U2 ( .A(n31), .B(n1), .Y(n34) );
  NAND2X2 U3 ( .A(n33), .B(n34), .Y(out6) );
  INVXLTH U4 ( .A(in6), .Y(n31) );
  INVXLTH U5 ( .A(n1), .Y(n32) );
  CLKNAND2X12 U6 ( .A(n37), .B(n38), .Y(n1) );
  XOR2X1 U7 ( .A(n46), .B(n1), .Y(out3) );
  XOR2X2 U9 ( .A(n44), .B(in2), .Y(n5) );
  CLKXOR2X4 U10 ( .A(n47), .B(n4), .Y(n3) );
  INVX2TH U11 ( .A(n2), .Y(n35) );
  NAND2X2 U12 ( .A(n2), .B(n3), .Y(n37) );
  INVX10 U13 ( .A(n3), .Y(n36) );
  XOR2XL U14 ( .A(in2), .B(n1), .Y(out2) );
  XOR2XL U15 ( .A(in5), .B(n1), .Y(out5) );
  INVXLTH U16 ( .A(n1), .Y(n40) );
  XOR2X1TH U17 ( .A(n47), .B(n1), .Y(out4) );
  CLKNAND2X8TH U18 ( .A(n35), .B(n36), .Y(n38) );
  XNOR2X4 U19 ( .A(in1), .B(n5), .Y(n2) );
  CLKNAND2X2TH U20 ( .A(n39), .B(n1), .Y(n42) );
  XOR2X4TH U22 ( .A(in6), .B(in5), .Y(n4) );
  INVXLTH U23 ( .A(in1), .Y(n39) );
  AND2X8 U8 ( .A(in1), .B(n40), .Y(n43) );
  CLKINVX40 U21 ( .A(n43), .Y(n41) );
  DLY1X1TH U24 ( .A(in3), .Y(n44) );
  INVXLTH U25 ( .A(n44), .Y(n45) );
  INVXLTH U26 ( .A(n45), .Y(n46) );
  DLY1X1TH U27 ( .A(in4), .Y(n47) );
  AND2X8 U28 ( .A(n41), .B(n42), .Y(n48) );
  CLKINVX40 U29 ( .A(n48), .Y(out1) );
endmodule


module all6_16 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n45, n46, n47, n48, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98;

  NAND3X2 U2 ( .A(n85), .B(n83), .C(n82), .Y(n26) );
  sign_xor_16 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR2XLTH U1 ( .A(n74), .B(n32), .Y(n45) );
  NOR2X8 U3 ( .A(n46), .B(n70), .Y(r3[0]) );
  INVX4 U4 ( .A(n45), .Y(n46) );
  INVX2TH U5 ( .A(n88), .Y(n74) );
  INVX1 U6 ( .A(n86), .Y(n70) );
  NOR2X3 U7 ( .A(n48), .B(n51), .Y(r4[0]) );
  INVXLTH U9 ( .A(n81), .Y(n64) );
  NAND3X2TH U10 ( .A(i5[1]), .B(i4[1]), .C(i6[1]), .Y(n31) );
  OR2XLTH U11 ( .A(n65), .B(n30), .Y(n47) );
  NOR3X1 U13 ( .A(n53), .B(n26), .C(n59), .Y(r5[2]) );
  NOR3X1 U14 ( .A(n51), .B(n28), .C(n60), .Y(r5[0]) );
  NOR2X2 U15 ( .A(n47), .B(n72), .Y(r2[2]) );
  NAND3X2 U16 ( .A(i5[2]), .B(n95), .C(i6[2]), .Y(n30) );
  NOR3X2 U17 ( .A(n29), .B(n71), .C(n63), .Y(r2[3]) );
  NOR3X1TH U18 ( .A(n58), .B(n25), .C(n62), .Y(r6[3]) );
  NOR2X3TH U19 ( .A(n50), .B(n66), .Y(r2[0]) );
  OR2XLTH U20 ( .A(n57), .B(n28), .Y(n48) );
  NAND3X2 U21 ( .A(n94), .B(n93), .C(n81), .Y(n27) );
  NOR3X1TH U22 ( .A(n55), .B(n26), .C(n59), .Y(r6[2]) );
  NAND3X4 U23 ( .A(n89), .B(n90), .C(n97), .Y(n32) );
  NOR3X4 U24 ( .A(n54), .B(n27), .C(n61), .Y(r5[1]) );
  NOR3X4 U25 ( .A(n31), .B(n69), .C(n64), .Y(r1[1]) );
  CLKINVX1 U26 ( .A(n94), .Y(n69) );
  CLKINVX1 U27 ( .A(n90), .Y(n51) );
  INVX1 U28 ( .A(n89), .Y(n57) );
  NOR3XL U29 ( .A(n30), .B(n68), .C(n65), .Y(r1[2]) );
  NOR3X4TH U30 ( .A(n29), .B(n71), .C(n67), .Y(r3[3]) );
  INVX2TH U31 ( .A(n87), .Y(n66) );
  OR2XLTH U33 ( .A(n74), .B(n32), .Y(n50) );
  NOR3X1TH U34 ( .A(n52), .B(n25), .C(n58), .Y(r4[3]) );
  NOR3X4 U35 ( .A(n57), .B(n28), .C(n60), .Y(r6[0]) );
  INVX2 U37 ( .A(n95), .Y(n59) );
  INVXLTH U38 ( .A(i4[3]), .Y(n62) );
  INVXLTH U40 ( .A(n77), .Y(n52) );
  NOR3X1TH U41 ( .A(n52), .B(n25), .C(n62), .Y(r5[3]) );
  INVXLTH U42 ( .A(n82), .Y(n65) );
  NOR3X4TH U43 ( .A(n30), .B(n72), .C(n68), .Y(r3[2]) );
  CLKINVX1TH U44 ( .A(i6[1]), .Y(n54) );
  CLKINVX1TH U45 ( .A(i5[1]), .Y(n56) );
  NOR3X4TH U46 ( .A(n54), .B(n27), .C(n56), .Y(r4[1]) );
  INVXLTH U47 ( .A(n79), .Y(n58) );
  INVXLTH U48 ( .A(n80), .Y(n71) );
  INVXLTH U49 ( .A(n78), .Y(n63) );
  NAND3X2TH U50 ( .A(i4[3]), .B(n79), .C(n77), .Y(n29) );
  INVXLTH U51 ( .A(n84), .Y(n67) );
  CLKINVX1TH U52 ( .A(i4[1]), .Y(n61) );
  INVXLTH U53 ( .A(n93), .Y(n73) );
  NOR3X1TH U54 ( .A(n29), .B(n67), .C(n63), .Y(r1[3]) );
  NOR3XLTH U56 ( .A(n53), .B(n26), .C(n55), .Y(r4[2]) );
  NOR3X4 U57 ( .A(n31), .B(n73), .C(n69), .Y(r3[1]) );
  CLKINVX1TH U58 ( .A(n97), .Y(n60) );
  INVXLTH U59 ( .A(i6[2]), .Y(n53) );
  INVXLTH U60 ( .A(n83), .Y(n72) );
  INVXLTH U61 ( .A(i5[2]), .Y(n55) );
  INVXLTH U62 ( .A(n85), .Y(n68) );
  AND3X8 U8 ( .A(n86), .B(n88), .C(n87), .Y(n75) );
  CLKINVX40 U12 ( .A(n75), .Y(n28) );
  AND3X8 U32 ( .A(n84), .B(n80), .C(n78), .Y(n76) );
  CLKINVX40 U36 ( .A(n76), .Y(n25) );
  DLY1X1TH U39 ( .A(i6[3]), .Y(n77) );
  DLY1X1TH U55 ( .A(i3[3]), .Y(n78) );
  DLY1X1TH U63 ( .A(i5[3]), .Y(n79) );
  DLY1X1TH U64 ( .A(i1[3]), .Y(n80) );
  DLY1X1TH U65 ( .A(i3[1]), .Y(n81) );
  DLY1X1TH U66 ( .A(i3[2]), .Y(n82) );
  DLY1X1TH U67 ( .A(i1[2]), .Y(n83) );
  DLY1X1TH U68 ( .A(i2[3]), .Y(n84) );
  DLY1X1TH U69 ( .A(i2[2]), .Y(n85) );
  DLY1X1TH U70 ( .A(i2[0]), .Y(n86) );
  DLY1X1TH U71 ( .A(i3[0]), .Y(n87) );
  DLY1X1TH U72 ( .A(i1[0]), .Y(n88) );
  DLY1X1TH U73 ( .A(i5[0]), .Y(n89) );
  DLY1X1TH U74 ( .A(i6[0]), .Y(n90) );
  DLY1X1TH U75 ( .A(n73), .Y(n91) );
  DLY1X1TH U76 ( .A(n64), .Y(n92) );
  DLY1X1TH U77 ( .A(i1[1]), .Y(n93) );
  DLY1X1TH U78 ( .A(i2[1]), .Y(n94) );
  DLY1X1TH U79 ( .A(i4[2]), .Y(n95) );
  NOR3BX4 U80 ( .AN(i5[1]), .B(n27), .C(n61), .Y(r6[1]) );
  NOR2BX8 U81 ( .AN(n96), .B(n31), .Y(r2[1]) );
  NOR2X8 U82 ( .A(n91), .B(n92), .Y(n96) );
  CLKBUFX40 U83 ( .A(i4[0]), .Y(n97) );
  OR3X8 U84 ( .A(n32), .B(n70), .C(n66), .Y(n98) );
  CLKINVX40 U85 ( .A(n98), .Y(r1[0]) );
endmodule


module sign_xor_15 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n4, n5, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39;

  CLKXOR2X12 U1 ( .A(n2), .B(n36), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(n33) );
  XOR2X1 U3 ( .A(in2), .B(n1), .Y(out2) );
  NAND2XLTH U4 ( .A(n32), .B(n1), .Y(n35) );
  XOR2X2 U5 ( .A(in6), .B(n1), .Y(out6) );
  XOR2XL U6 ( .A(in5), .B(n1), .Y(out5) );
  CLKNAND2X4 U7 ( .A(n30), .B(n31), .Y(out1) );
  NAND2XLTH U8 ( .A(n34), .B(n35), .Y(out3) );
  NAND2XLTH U9 ( .A(in1), .B(n29), .Y(n30) );
  NAND2XLTH U10 ( .A(n28), .B(n1), .Y(n31) );
  INVXLTH U11 ( .A(in1), .Y(n28) );
  INVXLTH U12 ( .A(n1), .Y(n29) );
  NAND2XL U13 ( .A(in3), .B(n33), .Y(n34) );
  INVXLTH U14 ( .A(in3), .Y(n32) );
  XOR2X3 U15 ( .A(in6), .B(in5), .Y(n4) );
  XNOR2X4 U16 ( .A(in1), .B(n5), .Y(n2) );
  XNOR2X4 U17 ( .A(n37), .B(n4), .Y(n36) );
  XOR2X2 U18 ( .A(in3), .B(in2), .Y(n5) );
  XOR2X1TH U19 ( .A(n39), .B(n1), .Y(out4) );
  DLY1X1TH U20 ( .A(in4), .Y(n37) );
  INVXLTH U21 ( .A(n37), .Y(n38) );
  INVXLTH U22 ( .A(n38), .Y(n39) );
endmodule


module all6_15 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85;

  NAND3X2 U1 ( .A(i1[3]), .B(n78), .C(n77), .Y(n25) );
  sign_xor_15 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X4 U2 ( .A(n32), .B(n69), .C(n62), .Y(r2[0]) );
  INVX2 U3 ( .A(n84), .Y(n69) );
  INVXL U4 ( .A(n82), .Y(n55) );
  NOR2X2 U5 ( .A(n45), .B(n61), .Y(r2[1]) );
  NOR3X4 U6 ( .A(n50), .B(n28), .C(n51), .Y(r4[0]) );
  OR2XLTH U7 ( .A(n70), .B(n31), .Y(n43) );
  CLKINVX1 U8 ( .A(n83), .Y(n62) );
  NOR2X2 U10 ( .A(n43), .B(n65), .Y(r3[1]) );
  NAND3X3 U11 ( .A(n80), .B(i4[1]), .C(i6[1]), .Y(n31) );
  INVX1 U12 ( .A(i1[1]), .Y(n70) );
  INVXL U13 ( .A(i2[1]), .Y(n65) );
  INVXLTH U14 ( .A(i3[1]), .Y(n61) );
  NOR3X4 U15 ( .A(n51), .B(n28), .C(n58), .Y(r6[0]) );
  NOR3X4 U16 ( .A(n32), .B(n69), .C(n66), .Y(r3[0]) );
  NAND3X4TH U17 ( .A(i2[1]), .B(i1[1]), .C(i3[1]), .Y(n27) );
  NOR2X2 U18 ( .A(n44), .B(n58), .Y(r5[0]) );
  NOR3X1 U20 ( .A(n30), .B(n67), .C(n59), .Y(r2[2]) );
  NOR3X2TH U21 ( .A(n47), .B(n26), .C(n52), .Y(r4[2]) );
  OR2X4 U22 ( .A(n50), .B(n28), .Y(n44) );
  NAND3X2 U23 ( .A(i5[0]), .B(i4[0]), .C(i6[0]), .Y(n32) );
  CLKINVX1 U24 ( .A(i2[0]), .Y(n66) );
  CLKINVX1TH U25 ( .A(i4[0]), .Y(n58) );
  CLKINVX1TH U26 ( .A(i5[0]), .Y(n51) );
  CLKINVX1TH U27 ( .A(i6[0]), .Y(n50) );
  NOR3X4TH U28 ( .A(n31), .B(n65), .C(n61), .Y(r1[1]) );
  NOR3X4TH U29 ( .A(n29), .B(n63), .C(n60), .Y(r1[3]) );
  NAND3X2TH U32 ( .A(i6[3]), .B(n76), .C(n75), .Y(n29) );
  NOR3X1TH U34 ( .A(n49), .B(n25), .C(n54), .Y(r4[3]) );
  NOR3X2TH U35 ( .A(n30), .B(n64), .C(n59), .Y(r1[2]) );
  OR2XLTH U36 ( .A(n31), .B(n70), .Y(n45) );
  OR2X1TH U37 ( .A(n53), .B(n56), .Y(n46) );
  NAND3X3 U38 ( .A(n81), .B(n82), .C(i6[2]), .Y(n30) );
  NOR3X1TH U39 ( .A(n49), .B(n25), .C(n57), .Y(r5[3]) );
  INVXLTH U40 ( .A(i1[3]), .Y(n68) );
  INVXLTH U41 ( .A(n80), .Y(n53) );
  INVXLTH U42 ( .A(n77), .Y(n60) );
  INVXLTH U43 ( .A(n78), .Y(n63) );
  NOR3X1TH U44 ( .A(n54), .B(n25), .C(n57), .Y(r6[3]) );
  NOR3X1TH U45 ( .A(n52), .B(n26), .C(n55), .Y(r6[2]) );
  NOR3X4TH U46 ( .A(n48), .B(n27), .C(n56), .Y(r5[1]) );
  INVX2 U48 ( .A(i2[2]), .Y(n64) );
  INVX2 U49 ( .A(n79), .Y(n59) );
  NOR3X1TH U50 ( .A(n29), .B(n68), .C(n63), .Y(r3[3]) );
  NOR3X1TH U51 ( .A(n29), .B(n68), .C(n60), .Y(r2[3]) );
  NOR3XLTH U52 ( .A(n30), .B(n67), .C(n64), .Y(r3[2]) );
  INVXLTH U53 ( .A(i4[1]), .Y(n56) );
  INVXLTH U54 ( .A(i6[1]), .Y(n48) );
  INVXLTH U55 ( .A(i6[2]), .Y(n47) );
  INVXLTH U56 ( .A(i6[3]), .Y(n49) );
  INVX2 U57 ( .A(i1[2]), .Y(n67) );
  INVXLTH U58 ( .A(n81), .Y(n52) );
  INVXLTH U59 ( .A(n75), .Y(n54) );
  INVXLTH U60 ( .A(n76), .Y(n57) );
  NAND2BX8 U9 ( .AN(n46), .B(n72), .Y(n71) );
  CLKINVX40 U19 ( .A(n71), .Y(r6[1]) );
  CLKINVX40 U30 ( .A(n27), .Y(n72) );
  AND3X8 U31 ( .A(n84), .B(n83), .C(i2[0]), .Y(n73) );
  CLKINVX40 U33 ( .A(n73), .Y(n28) );
  AND3X8 U47 ( .A(i2[2]), .B(i1[2]), .C(n79), .Y(n74) );
  CLKINVX40 U61 ( .A(n74), .Y(n26) );
  NOR3BX4 U62 ( .AN(i6[2]), .B(n26), .C(n55), .Y(r5[2]) );
  NOR3BX4 U63 ( .AN(i6[1]), .B(n27), .C(n53), .Y(r4[1]) );
  DLY1X1TH U64 ( .A(i5[3]), .Y(n75) );
  DLY1X1TH U65 ( .A(i4[3]), .Y(n76) );
  DLY1X1TH U66 ( .A(i3[3]), .Y(n77) );
  DLY1X1TH U67 ( .A(i2[3]), .Y(n78) );
  DLY1X1TH U68 ( .A(i3[2]), .Y(n79) );
  DLY1X1TH U69 ( .A(i5[1]), .Y(n80) );
  DLY1X1TH U70 ( .A(i5[2]), .Y(n81) );
  DLY1X1TH U71 ( .A(i4[2]), .Y(n82) );
  DLY1X1TH U72 ( .A(i3[0]), .Y(n83) );
  DLY1X1TH U73 ( .A(i1[0]), .Y(n84) );
  OR3X8 U74 ( .A(n32), .B(n66), .C(n62), .Y(n85) );
  CLKINVX40 U75 ( .A(n85), .Y(r1[0]) );
endmodule


module sign_xor_14 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n4, n5, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39;

  NAND2XL U1 ( .A(in3), .B(n24), .Y(n25) );
  INVXL U2 ( .A(n1), .Y(n24) );
  CLKNAND2X4 U3 ( .A(n28), .B(n29), .Y(out5) );
  XOR2X3 U4 ( .A(in6), .B(in5), .Y(n4) );
  XOR2X1 U5 ( .A(in4), .B(n1), .Y(out4) );
  NAND2X8 U6 ( .A(n32), .B(n33), .Y(n1) );
  NAND2X2 U7 ( .A(n2), .B(n31), .Y(n32) );
  INVX2 U8 ( .A(n34), .Y(n31) );
  NAND2X2 U9 ( .A(n25), .B(n26), .Y(out3) );
  NAND2X3 U10 ( .A(n34), .B(n30), .Y(n33) );
  NAND2XLTH U11 ( .A(n23), .B(n1), .Y(n26) );
  INVXLTH U12 ( .A(in3), .Y(n23) );
  INVX10TH U13 ( .A(n2), .Y(n30) );
  XOR2X3TH U16 ( .A(in3), .B(in2), .Y(n5) );
  NAND2XLTH U18 ( .A(n27), .B(n1), .Y(n29) );
  INVXLTH U19 ( .A(in5), .Y(n27) );
  XNOR2X4 U21 ( .A(n38), .B(n5), .Y(n2) );
  XNOR2X4 U22 ( .A(in4), .B(n4), .Y(n34) );
  XNOR2X1 U14 ( .A(n39), .B(n1), .Y(out1) );
  XNOR2X1 U15 ( .A(n35), .B(n1), .Y(out2) );
  CLKINVX40 U17 ( .A(in2), .Y(n35) );
  AND2X8 U20 ( .A(in5), .B(n24), .Y(n36) );
  CLKINVX40 U23 ( .A(n36), .Y(n28) );
  XNOR2X1 U24 ( .A(n37), .B(n1), .Y(out6) );
  CLKINVX40 U25 ( .A(in6), .Y(n37) );
  DLY1X1TH U26 ( .A(in1), .Y(n38) );
  INVXLTH U27 ( .A(n38), .Y(n39) );
endmodule


module all6_14 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82;

  NAND3X2 U2 ( .A(i2[2]), .B(i1[2]), .C(i3[2]), .Y(n26) );
  NOR3X1 U34 ( .A(n55), .B(n26), .C(n59), .Y(r6[2]) );
  sign_xor_14 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X1 U1 ( .A(n30), .B(n73), .C(n69), .Y(r3[2]) );
  OR2X4 U3 ( .A(n58), .B(n54), .Y(n50) );
  INVXL U4 ( .A(n79), .Y(n52) );
  INVXL U5 ( .A(i3[2]), .Y(n66) );
  NOR3X1TH U6 ( .A(n29), .B(n72), .C(n67), .Y(r3[3]) );
  NOR3X4TH U7 ( .A(n32), .B(n70), .C(n65), .Y(r1[0]) );
  INVX2 U8 ( .A(n81), .Y(n65) );
  NOR3X1 U9 ( .A(n57), .B(n25), .C(n61), .Y(r6[3]) );
  NOR3XL U10 ( .A(n30), .B(n73), .C(n66), .Y(r2[2]) );
  CLKINVX1TH U11 ( .A(i4[0]), .Y(n60) );
  INVXLTH U12 ( .A(i5[1]), .Y(n56) );
  NAND3X3TH U13 ( .A(i5[1]), .B(i4[1]), .C(i6[1]), .Y(n31) );
  INVX2TH U14 ( .A(i5[0]), .Y(n58) );
  NAND3X3 U15 ( .A(n81), .B(i1[0]), .C(i2[0]), .Y(n28) );
  NOR3X4TH U16 ( .A(n52), .B(n26), .C(n55), .Y(r4[2]) );
  NOR3X4TH U17 ( .A(n32), .B(n74), .C(n70), .Y(r3[0]) );
  NOR3X1TH U18 ( .A(n29), .B(n72), .C(n63), .Y(r2[3]) );
  NOR3X2 U19 ( .A(n31), .B(n71), .C(n64), .Y(r2[1]) );
  NOR3X4TH U20 ( .A(n53), .B(n27), .C(n56), .Y(r4[1]) );
  INVX1TH U23 ( .A(i1[0]), .Y(n74) );
  NAND3X4TH U24 ( .A(i5[0]), .B(i4[0]), .C(i6[0]), .Y(n32) );
  NAND3X4TH U25 ( .A(n79), .B(n80), .C(i5[2]), .Y(n30) );
  NOR3X1TH U26 ( .A(n51), .B(n25), .C(n57), .Y(r4[3]) );
  NOR2X2TH U27 ( .A(n50), .B(n28), .Y(r4[0]) );
  INVXLTH U28 ( .A(i2[3]), .Y(n67) );
  INVXLTH U29 ( .A(n77), .Y(n57) );
  INVXLTH U30 ( .A(n76), .Y(n51) );
  NAND3X2TH U31 ( .A(i2[3]), .B(n78), .C(n75), .Y(n25) );
  INVXLTH U32 ( .A(i4[3]), .Y(n61) );
  INVXLTH U33 ( .A(i4[1]), .Y(n62) );
  INVXLTH U35 ( .A(n78), .Y(n72) );
  NAND3X2TH U36 ( .A(i4[3]), .B(n77), .C(n76), .Y(n29) );
  INVXLTH U37 ( .A(n75), .Y(n63) );
  INVXLTH U38 ( .A(i1[2]), .Y(n73) );
  CLKINVX1TH U39 ( .A(i2[1]), .Y(n68) );
  NOR3X1TH U40 ( .A(n29), .B(n67), .C(n63), .Y(r1[3]) );
  CLKINVX1TH U41 ( .A(i2[0]), .Y(n70) );
  NOR3X1TH U42 ( .A(n51), .B(n25), .C(n61), .Y(r5[3]) );
  NOR3X1TH U43 ( .A(n53), .B(n27), .C(n62), .Y(r5[1]) );
  NOR3X4TH U44 ( .A(n31), .B(n71), .C(n68), .Y(r3[1]) );
  NAND3X2TH U45 ( .A(i2[1]), .B(i1[1]), .C(i3[1]), .Y(n27) );
  NOR3X4TH U46 ( .A(n31), .B(n68), .C(n64), .Y(r1[1]) );
  NOR3X4TH U47 ( .A(n32), .B(n74), .C(n65), .Y(r2[0]) );
  INVXLTH U49 ( .A(i6[0]), .Y(n54) );
  INVXLTH U50 ( .A(i1[1]), .Y(n71) );
  INVX2 U51 ( .A(i2[2]), .Y(n69) );
  NOR3XLTH U52 ( .A(n30), .B(n69), .C(n66), .Y(r1[2]) );
  INVXLTH U54 ( .A(i6[1]), .Y(n53) );
  INVXLTH U55 ( .A(i5[2]), .Y(n55) );
  INVXLTH U56 ( .A(n80), .Y(n59) );
  INVXLTH U57 ( .A(i3[1]), .Y(n64) );
  NOR3BX4 U21 ( .AN(i6[0]), .B(n28), .C(n60), .Y(r5[0]) );
  NOR3BX4 U22 ( .AN(n79), .B(n26), .C(n59), .Y(r5[2]) );
  DLY1X1TH U48 ( .A(i3[3]), .Y(n75) );
  DLY1X1TH U53 ( .A(i6[3]), .Y(n76) );
  DLY1X1TH U58 ( .A(i5[3]), .Y(n77) );
  DLY1X1TH U59 ( .A(i1[3]), .Y(n78) );
  DLY1X1TH U60 ( .A(i6[2]), .Y(n79) );
  DLY1X1TH U61 ( .A(i4[2]), .Y(n80) );
  DLY1X1TH U62 ( .A(i3[0]), .Y(n81) );
  NOR3BX4 U63 ( .AN(i5[1]), .B(n27), .C(n62), .Y(r6[1]) );
  OR3X8 U64 ( .A(n58), .B(n28), .C(n60), .Y(n82) );
  CLKINVX40 U65 ( .A(n82), .Y(r6[0]) );
endmodule


module sign_xor_13 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n3, n4, n5, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42;

  XOR2X1 U1 ( .A(in6), .B(n1), .Y(out6) );
  CLKXOR2X12 U2 ( .A(n39), .B(n3), .Y(n1) );
  NAND2XLTH U3 ( .A(in3), .B(n32), .Y(n33) );
  NAND2XLTH U4 ( .A(n31), .B(n1), .Y(n34) );
  NAND2X2 U5 ( .A(n33), .B(n34), .Y(out3) );
  INVXLTH U6 ( .A(in3), .Y(n31) );
  INVXL U7 ( .A(n1), .Y(n32) );
  CLKXOR2X2TH U8 ( .A(in4), .B(n4), .Y(n3) );
  CLKXOR2X2TH U9 ( .A(in2), .B(n1), .Y(out2) );
  CLKNAND2X2TH U10 ( .A(n37), .B(n38), .Y(out4) );
  XOR2XLTH U11 ( .A(in5), .B(n1), .Y(out5) );
  XOR2X4 U12 ( .A(in6), .B(in5), .Y(n4) );
  INVX1TH U13 ( .A(n1), .Y(n36) );
  NAND2X1TH U14 ( .A(in4), .B(n36), .Y(n37) );
  NAND2XLTH U15 ( .A(n35), .B(n1), .Y(n38) );
  INVXLTH U16 ( .A(in4), .Y(n35) );
  XOR2X1TH U17 ( .A(n42), .B(n1), .Y(out1) );
  XOR2X2 U18 ( .A(n40), .B(n5), .Y(n39) );
  XOR2X3TH U19 ( .A(in3), .B(in2), .Y(n5) );
  DLY1X1TH U20 ( .A(in1), .Y(n40) );
  INVXLTH U21 ( .A(n40), .Y(n41) );
  INVXLTH U22 ( .A(n41), .Y(n42) );
endmodule


module all6_13 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80;

  NOR3X1 U50 ( .A(n30), .B(n66), .C(n57), .Y(r2[2]) );
  sign_xor_13 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NAND3X2 U1 ( .A(i6[3]), .B(n74), .C(n72), .Y(n29) );
  NAND3X2 U2 ( .A(i3[2]), .B(n75), .C(n73), .Y(n26) );
  NAND3X2 U3 ( .A(i5[1]), .B(i4[1]), .C(i6[1]), .Y(n31) );
  CLKINVX2TH U4 ( .A(n76), .Y(n63) );
  CLKNAND2X2 U5 ( .A(i4[0]), .B(i6[0]), .Y(n37) );
  NAND2X4 U6 ( .A(n78), .B(n38), .Y(n32) );
  INVX4 U7 ( .A(n37), .Y(n38) );
  NOR3X4 U8 ( .A(n32), .B(n67), .C(n64), .Y(r3[0]) );
  NOR2X4 U10 ( .A(n57), .B(n62), .Y(n39) );
  NOR2XLTH U11 ( .A(n40), .B(n30), .Y(r1[2]) );
  INVX2 U12 ( .A(n39), .Y(n40) );
  NAND3X3 U13 ( .A(n77), .B(i5[2]), .C(n79), .Y(n30) );
  NAND3X2 U15 ( .A(i2[0]), .B(i1[0]), .C(i3[0]), .Y(n28) );
  NOR3X1TH U16 ( .A(n45), .B(n25), .C(n49), .Y(r4[3]) );
  NOR3X1TH U17 ( .A(n29), .B(n65), .C(n58), .Y(r2[3]) );
  NOR2X2 U18 ( .A(n41), .B(n28), .Y(r4[0]) );
  OR2XLTH U19 ( .A(n48), .B(n52), .Y(n41) );
  NOR2X2 U20 ( .A(n44), .B(n27), .Y(r6[1]) );
  OR2X2 U21 ( .A(n55), .B(n51), .Y(n44) );
  INVX2 U22 ( .A(n78), .Y(n52) );
  NOR2X3 U23 ( .A(n43), .B(n48), .Y(r5[0]) );
  INVX1 U24 ( .A(i5[2]), .Y(n50) );
  CLKINVX1 U25 ( .A(i3[0]), .Y(n59) );
  NAND3X2 U26 ( .A(i3[1]), .B(i1[1]), .C(n76), .Y(n27) );
  CLKINVX1TH U27 ( .A(i2[0]), .Y(n64) );
  NOR3X4 U28 ( .A(n31), .B(n68), .C(n60), .Y(r2[1]) );
  INVXL U29 ( .A(i1[1]), .Y(n68) );
  NOR3X4 U30 ( .A(n46), .B(n26), .C(n50), .Y(r4[2]) );
  NOR3X1TH U31 ( .A(n45), .B(n25), .C(n53), .Y(r5[3]) );
  INVXLTH U32 ( .A(n77), .Y(n54) );
  INVXLTH U33 ( .A(i4[0]), .Y(n56) );
  NOR3X4TH U34 ( .A(n29), .B(n65), .C(n61), .Y(r3[3]) );
  OR2XLTH U35 ( .A(n50), .B(n54), .Y(n42) );
  OR2XLTH U36 ( .A(n56), .B(n28), .Y(n43) );
  NOR2XLTH U37 ( .A(n42), .B(n26), .Y(r6[2]) );
  INVXLTH U38 ( .A(n71), .Y(n65) );
  INVXLTH U39 ( .A(i4[1]), .Y(n55) );
  INVXLTH U40 ( .A(i6[1]), .Y(n47) );
  INVXLTH U41 ( .A(i5[1]), .Y(n51) );
  CLKINVX1TH U42 ( .A(i6[0]), .Y(n48) );
  CLKINVX1TH U43 ( .A(i1[0]), .Y(n67) );
  NOR3X1TH U44 ( .A(n29), .B(n61), .C(n58), .Y(r1[3]) );
  NOR3X1TH U45 ( .A(n30), .B(n66), .C(n62), .Y(r3[2]) );
  NOR3X2 U46 ( .A(n31), .B(n68), .C(n63), .Y(r3[1]) );
  INVXLTH U47 ( .A(i3[3]), .Y(n58) );
  INVXLTH U48 ( .A(n70), .Y(n61) );
  INVXLTH U49 ( .A(n72), .Y(n49) );
  INVXLTH U51 ( .A(n74), .Y(n53) );
  NAND3X2TH U52 ( .A(i3[3]), .B(n71), .C(n70), .Y(n25) );
  INVXLTH U53 ( .A(i6[3]), .Y(n45) );
  INVXLTH U54 ( .A(i3[1]), .Y(n60) );
  NOR3X1TH U55 ( .A(n52), .B(n28), .C(n56), .Y(r6[0]) );
  NOR3X1TH U56 ( .A(n49), .B(n25), .C(n53), .Y(r6[3]) );
  NOR3X4TH U57 ( .A(n47), .B(n27), .C(n55), .Y(r5[1]) );
  NOR3X2 U58 ( .A(n31), .B(n63), .C(n60), .Y(r1[1]) );
  NOR3X2 U59 ( .A(n47), .B(n27), .C(n51), .Y(r4[1]) );
  INVXLTH U61 ( .A(n75), .Y(n66) );
  INVXLTH U62 ( .A(n73), .Y(n62) );
  INVXLTH U63 ( .A(n79), .Y(n46) );
  INVXLTH U64 ( .A(i3[2]), .Y(n57) );
  OR3X8 U9 ( .A(n32), .B(n67), .C(n59), .Y(n69) );
  CLKINVX40 U14 ( .A(n69), .Y(r2[0]) );
  NOR3BX4 U60 ( .AN(n79), .B(n26), .C(n54), .Y(r5[2]) );
  DLY1X1TH U65 ( .A(i2[3]), .Y(n70) );
  DLY1X1TH U66 ( .A(i1[3]), .Y(n71) );
  DLY1X1TH U67 ( .A(i5[3]), .Y(n72) );
  DLY1X1TH U68 ( .A(i2[2]), .Y(n73) );
  DLY1X1TH U69 ( .A(i4[3]), .Y(n74) );
  DLY1X1TH U70 ( .A(i1[2]), .Y(n75) );
  DLY1X1TH U71 ( .A(i2[1]), .Y(n76) );
  DLY1X1TH U72 ( .A(i4[2]), .Y(n77) );
  DLY1X1TH U73 ( .A(i5[0]), .Y(n78) );
  DLY1X1TH U74 ( .A(i6[2]), .Y(n79) );
  NOR3BX4 U75 ( .AN(n80), .B(n64), .C(n59), .Y(r1[0]) );
  CLKINVX40 U76 ( .A(n32), .Y(n80) );
endmodule


module sign_xor_12 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44;

  NAND2X5 U1 ( .A(n40), .B(n41), .Y(n1) );
  XNOR2X4 U2 ( .A(in1), .B(n5), .Y(n2) );
  NAND2X2 U3 ( .A(n36), .B(n37), .Y(out1) );
  BUFX8 U4 ( .A(in6), .Y(n26) );
  BUFX6 U5 ( .A(in5), .Y(n27) );
  BUFX6 U6 ( .A(in3), .Y(n28) );
  BUFX8 U7 ( .A(in2), .Y(n29) );
  XOR2X8 U8 ( .A(in4), .B(n4), .Y(n3) );
  XOR2X1 U9 ( .A(in4), .B(n1), .Y(out4) );
  XOR2X4 U10 ( .A(n28), .B(n29), .Y(n5) );
  NAND2XLTH U11 ( .A(n29), .B(n31), .Y(n32) );
  NAND2X1 U12 ( .A(n30), .B(n1), .Y(n33) );
  CLKNAND2X4 U13 ( .A(n32), .B(n33), .Y(out2) );
  INVXLTH U14 ( .A(n29), .Y(n30) );
  INVX4 U15 ( .A(n1), .Y(n31) );
  INVX3 U16 ( .A(n2), .Y(n38) );
  CLKNAND2X2TH U17 ( .A(n43), .B(n44), .Y(out6) );
  XOR2X2 U18 ( .A(n28), .B(n1), .Y(out3) );
  CLKINVX2 U19 ( .A(n1), .Y(n35) );
  XOR2X4 U20 ( .A(n26), .B(n27), .Y(n4) );
  NAND2X2TH U21 ( .A(in1), .B(n35), .Y(n36) );
  NAND2XL U22 ( .A(n34), .B(n1), .Y(n37) );
  INVXLTH U23 ( .A(in1), .Y(n34) );
  XOR2XLTH U24 ( .A(n27), .B(n1), .Y(out5) );
  NAND2XLTH U25 ( .A(n42), .B(n1), .Y(n44) );
  CLKNAND2X4 U26 ( .A(n38), .B(n39), .Y(n41) );
  INVX2TH U27 ( .A(n3), .Y(n39) );
  NAND2X4 U28 ( .A(n2), .B(n3), .Y(n40) );
  NAND2X1 U29 ( .A(n26), .B(n35), .Y(n43) );
  INVXLTH U30 ( .A(n26), .Y(n42) );
endmodule


module all6_12 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95;

  NAND3X2 U5 ( .A(i5[3]), .B(i4[3]), .C(i6[3]), .Y(n29) );
  sign_xor_12 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NAND3X3 U1 ( .A(n89), .B(n90), .C(i4[1]), .Y(n31) );
  INVX2 U2 ( .A(n88), .Y(n71) );
  NOR3X2 U3 ( .A(n30), .B(n78), .C(n69), .Y(r2[2]) );
  NOR3X4 U4 ( .A(n30), .B(n78), .C(n74), .Y(r3[2]) );
  NAND3X2 U6 ( .A(i5[2]), .B(i4[2]), .C(n85), .Y(n30) );
  NOR2X2 U7 ( .A(n54), .B(n72), .Y(r1[0]) );
  NOR3X2 U8 ( .A(n30), .B(n74), .C(n69), .Y(r1[2]) );
  NOR3X2 U9 ( .A(n60), .B(n28), .C(n64), .Y(r4[0]) );
  INVX2TH U11 ( .A(i1[0]), .Y(n55) );
  NOR3X1TH U12 ( .A(n61), .B(n25), .C(n65), .Y(r6[3]) );
  OR2X2 U13 ( .A(n55), .B(n56), .Y(n28) );
  NOR2X4 U15 ( .A(n52), .B(n64), .Y(r6[0]) );
  INVX2TH U16 ( .A(i4[2]), .Y(n66) );
  INVXLTH U17 ( .A(i4[0]), .Y(n68) );
  INVXLTH U18 ( .A(i5[2]), .Y(n62) );
  NAND3X4TH U19 ( .A(n91), .B(n92), .C(i4[0]), .Y(n32) );
  OR2XLTH U20 ( .A(n62), .B(n66), .Y(n51) );
  OR2X2TH U21 ( .A(n68), .B(n28), .Y(n52) );
  NOR3X4 U22 ( .A(n32), .B(n55), .C(n76), .Y(r3[0]) );
  NOR2XLTH U23 ( .A(n51), .B(n26), .Y(r6[2]) );
  NAND3X2 U24 ( .A(n87), .B(n86), .C(n84), .Y(n26) );
  NOR3X1TH U25 ( .A(n58), .B(n26), .C(n62), .Y(r4[2]) );
  NOR3X2TH U26 ( .A(n29), .B(n77), .C(n73), .Y(r3[3]) );
  INVXLTH U27 ( .A(n85), .Y(n58) );
  INVXLTH U28 ( .A(n89), .Y(n63) );
  INVXLTH U29 ( .A(n90), .Y(n59) );
  INVXLTH U30 ( .A(n86), .Y(n78) );
  INVXLTH U31 ( .A(n84), .Y(n69) );
  INVXLTH U32 ( .A(i2[3]), .Y(n73) );
  NAND2XLTH U33 ( .A(i3[0]), .B(i2[0]), .Y(n56) );
  INVXLTH U34 ( .A(i2[0]), .Y(n76) );
  CLKINVX1TH U35 ( .A(i3[0]), .Y(n72) );
  NOR3X4 U36 ( .A(n60), .B(n28), .C(n68), .Y(r5[0]) );
  OR2XLTH U37 ( .A(n59), .B(n63), .Y(n53) );
  OR2XLTH U38 ( .A(n32), .B(n76), .Y(n54) );
  NOR3X2 U39 ( .A(n29), .B(n73), .C(n70), .Y(r1[3]) );
  NOR3X1TH U40 ( .A(n58), .B(n26), .C(n66), .Y(r5[2]) );
  NOR3X2 U42 ( .A(n59), .B(n27), .C(n67), .Y(r5[1]) );
  NOR3X1TH U43 ( .A(n57), .B(n25), .C(n61), .Y(r4[3]) );
  INVXLTH U44 ( .A(n93), .Y(n77) );
  NOR3X4TH U45 ( .A(n31), .B(n79), .C(n75), .Y(r3[1]) );
  NOR3X1TH U46 ( .A(n29), .B(n77), .C(n70), .Y(r2[3]) );
  INVXLTH U47 ( .A(i6[3]), .Y(n57) );
  INVXLTH U48 ( .A(i4[3]), .Y(n65) );
  INVXLTH U49 ( .A(i5[3]), .Y(n61) );
  NAND3X2TH U50 ( .A(i2[3]), .B(n93), .C(i3[3]), .Y(n25) );
  INVXLTH U51 ( .A(i4[1]), .Y(n67) );
  NOR3X1TH U52 ( .A(n57), .B(n25), .C(n65), .Y(r5[3]) );
  INVXLTH U53 ( .A(i1[1]), .Y(n79) );
  INVXLTH U54 ( .A(n94), .Y(n75) );
  INVXLTH U55 ( .A(i3[3]), .Y(n70) );
  INVXLTH U56 ( .A(n92), .Y(n60) );
  INVXLTH U57 ( .A(n91), .Y(n64) );
  NOR3X4TH U58 ( .A(n32), .B(n55), .C(n72), .Y(r2[0]) );
  NOR3X2 U59 ( .A(n31), .B(n75), .C(n71), .Y(r1[1]) );
  INVXLTH U61 ( .A(n87), .Y(n74) );
  AND3X8 U10 ( .A(n94), .B(i1[1]), .C(n88), .Y(n80) );
  CLKINVX40 U14 ( .A(n80), .Y(n27) );
  NAND3BX4 U41 ( .AN(n63), .B(n80), .C(i4[1]), .Y(n81) );
  CLKINVX40 U60 ( .A(n81), .Y(r6[1]) );
  NAND3BX4 U62 ( .AN(n31), .B(i1[1]), .C(n83), .Y(n82) );
  CLKINVX40 U63 ( .A(n82), .Y(r2[1]) );
  CLKINVX40 U64 ( .A(n71), .Y(n83) );
  DLY1X1TH U65 ( .A(i3[2]), .Y(n84) );
  DLY1X1TH U66 ( .A(i6[2]), .Y(n85) );
  DLY1X1TH U67 ( .A(i1[2]), .Y(n86) );
  DLY1X1TH U68 ( .A(i2[2]), .Y(n87) );
  DLY1X1TH U69 ( .A(i3[1]), .Y(n88) );
  DLY1X1TH U70 ( .A(i5[1]), .Y(n89) );
  DLY1X1TH U71 ( .A(i6[1]), .Y(n90) );
  DLY1X1TH U72 ( .A(i5[0]), .Y(n91) );
  DLY1X1TH U73 ( .A(i6[0]), .Y(n92) );
  DLY1X1TH U74 ( .A(i1[3]), .Y(n93) );
  DLY1X1TH U75 ( .A(i2[1]), .Y(n94) );
  OR2X8 U76 ( .A(n53), .B(n27), .Y(n95) );
  CLKINVX40 U77 ( .A(n95), .Y(r4[1]) );
endmodule


module sign_xor_11 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n4, n5, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37;

  NAND2X6 U1 ( .A(in6), .B(n23), .Y(n24) );
  NAND2X4 U2 ( .A(n22), .B(in5), .Y(n25) );
  CLKNAND2X8 U3 ( .A(n24), .B(n25), .Y(n4) );
  INVXLTH U4 ( .A(in6), .Y(n22) );
  INVX5 U5 ( .A(in5), .Y(n23) );
  NAND2X4 U6 ( .A(in3), .B(n27), .Y(n28) );
  NAND2X6 U7 ( .A(n26), .B(in2), .Y(n29) );
  CLKNAND2X8 U8 ( .A(n28), .B(n29), .Y(n5) );
  INVX2 U9 ( .A(in3), .Y(n26) );
  CLKINVX1 U10 ( .A(in2), .Y(n27) );
  XNOR2X2 U11 ( .A(in1), .B(n5), .Y(n2) );
  XOR2X1 U12 ( .A(in6), .B(n1), .Y(out6) );
  CLKNAND2X2TH U13 ( .A(n32), .B(n33), .Y(out1) );
  NAND2X1TH U14 ( .A(in1), .B(n31), .Y(n32) );
  XOR2X1 U15 ( .A(in2), .B(n1), .Y(out2) );
  NAND2XL U16 ( .A(n30), .B(n1), .Y(n33) );
  INVXLTH U17 ( .A(in1), .Y(n30) );
  INVXL U18 ( .A(n1), .Y(n31) );
  XOR2XL U19 ( .A(n37), .B(n1), .Y(out4) );
  XOR2X1 U20 ( .A(in3), .B(n1), .Y(out3) );
  XOR2X8 U21 ( .A(n2), .B(n34), .Y(n1) );
  XOR2XLTH U22 ( .A(in5), .B(n1), .Y(out5) );
  XNOR2X4 U23 ( .A(n35), .B(n4), .Y(n34) );
  DLY1X1TH U24 ( .A(in4), .Y(n35) );
  INVXLTH U25 ( .A(n35), .Y(n36) );
  INVXLTH U26 ( .A(n36), .Y(n37) );
endmodule


module all6_11 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n44, n45, n46, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87;

  sign_xor_11 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X1 U1 ( .A(n30), .B(n69), .C(n61), .Y(r2[2]) );
  AND2XLTH U3 ( .A(n72), .B(i6[1]), .Y(n44) );
  NAND2X2 U4 ( .A(i5[1]), .B(n44), .Y(n31) );
  NOR2X2 U5 ( .A(n45), .B(n31), .Y(r3[1]) );
  NOR3XLTH U7 ( .A(n50), .B(n26), .C(n57), .Y(r5[2]) );
  NOR3X2 U8 ( .A(n31), .B(n65), .C(n60), .Y(r1[1]) );
  NOR3X1TH U9 ( .A(n30), .B(n64), .C(n61), .Y(r1[2]) );
  INVX2 U10 ( .A(i1[1]), .Y(n68) );
  INVX1TH U11 ( .A(i2[1]), .Y(n65) );
  NAND3X2TH U12 ( .A(i2[3]), .B(n74), .C(n73), .Y(n25) );
  NOR3X2TH U13 ( .A(n53), .B(n26), .C(n57), .Y(r6[2]) );
  INVXLTH U14 ( .A(i5[2]), .Y(n53) );
  NOR3X1 U17 ( .A(n49), .B(n27), .C(n52), .Y(r4[1]) );
  OR2XLTH U18 ( .A(n68), .B(n65), .Y(n45) );
  INVXLTH U20 ( .A(n75), .Y(n55) );
  NOR3X1TH U21 ( .A(n51), .B(n25), .C(n55), .Y(r6[3]) );
  NOR3X1TH U22 ( .A(n29), .B(n67), .C(n59), .Y(r2[3]) );
  INVXLTH U23 ( .A(i5[3]), .Y(n51) );
  INVX2TH U24 ( .A(i6[2]), .Y(n50) );
  NOR3X1TH U25 ( .A(n32), .B(n66), .C(n62), .Y(r1[0]) );
  OR2XLTH U26 ( .A(n49), .B(n56), .Y(n46) );
  NOR3X1TH U29 ( .A(n50), .B(n26), .C(n53), .Y(r4[2]) );
  NOR3X4 U30 ( .A(n54), .B(n28), .C(n58), .Y(r6[0]) );
  NOR3X1TH U31 ( .A(n30), .B(n69), .C(n64), .Y(r3[2]) );
  INVXLTH U32 ( .A(i6[3]), .Y(n48) );
  INVXLTH U33 ( .A(n74), .Y(n67) );
  INVXLTH U34 ( .A(n72), .Y(n56) );
  NOR3X1TH U35 ( .A(n48), .B(n25), .C(n55), .Y(r5[3]) );
  CLKINVX1TH U36 ( .A(i4[0]), .Y(n58) );
  INVXLTH U37 ( .A(i6[1]), .Y(n49) );
  NOR3X1TH U39 ( .A(n29), .B(n67), .C(n63), .Y(r3[3]) );
  INVXLTH U40 ( .A(i3[1]), .Y(n60) );
  NAND3X2TH U41 ( .A(i5[3]), .B(n75), .C(i6[3]), .Y(n29) );
  INVXLTH U42 ( .A(i2[3]), .Y(n63) );
  INVXLTH U43 ( .A(n73), .Y(n59) );
  INVXLTH U44 ( .A(i2[0]), .Y(n66) );
  NOR3X4TH U45 ( .A(n52), .B(n27), .C(n56), .Y(r6[1]) );
  INVXLTH U46 ( .A(i3[0]), .Y(n62) );
  NAND3X3TH U47 ( .A(n87), .B(i4[0]), .C(i6[0]), .Y(n32) );
  CLKINVX1TH U48 ( .A(i1[0]), .Y(n70) );
  NOR3X1TH U49 ( .A(n29), .B(n63), .C(n59), .Y(r1[3]) );
  NOR3X4TH U50 ( .A(n32), .B(n70), .C(n62), .Y(r2[0]) );
  NOR3X4TH U51 ( .A(n32), .B(n70), .C(n66), .Y(r3[0]) );
  INVXLTH U53 ( .A(i5[1]), .Y(n52) );
  INVXLTH U55 ( .A(n80), .Y(n69) );
  INVXLTH U56 ( .A(n76), .Y(n64) );
  INVXLTH U57 ( .A(n78), .Y(n57) );
  INVXLTH U58 ( .A(n77), .Y(n61) );
  CLKINVX1TH U59 ( .A(n87), .Y(n54) );
  AND3X8 U2 ( .A(i2[0]), .B(i1[0]), .C(i3[0]), .Y(n71) );
  CLKINVX40 U6 ( .A(n71), .Y(n28) );
  NOR3BX4 U15 ( .AN(i6[0]), .B(n28), .C(n58), .Y(r5[0]) );
  AND3X8 U16 ( .A(i6[0]), .B(n71), .C(n87), .Y(r4[0]) );
  DLY1X1TH U19 ( .A(i4[1]), .Y(n72) );
  DLY1X1TH U27 ( .A(i3[3]), .Y(n73) );
  DLY1X1TH U28 ( .A(i1[3]), .Y(n74) );
  DLY1X1TH U38 ( .A(i4[3]), .Y(n75) );
  DLY1X1TH U52 ( .A(i2[2]), .Y(n76) );
  DLY1X1TH U54 ( .A(i3[2]), .Y(n77) );
  DLY1X1TH U60 ( .A(i4[2]), .Y(n78) );
  INVXLTH U61 ( .A(n50), .Y(n79) );
  CLKBUFX40 U62 ( .A(i1[2]), .Y(n80) );
  AND3X8 U63 ( .A(i2[1]), .B(i1[1]), .C(i3[1]), .Y(n81) );
  CLKINVX40 U64 ( .A(n81), .Y(n27) );
  AND3X8 U65 ( .A(i5[2]), .B(n78), .C(n79), .Y(n82) );
  CLKINVX40 U66 ( .A(n82), .Y(n30) );
  AND3X8 U67 ( .A(n76), .B(n80), .C(n77), .Y(n83) );
  CLKINVX40 U68 ( .A(n83), .Y(n26) );
  NAND3BX4 U69 ( .AN(n31), .B(n85), .C(i3[1]), .Y(n84) );
  CLKINVX40 U70 ( .A(n84), .Y(r2[1]) );
  CLKINVX40 U71 ( .A(n68), .Y(n85) );
  NOR3BX4 U72 ( .AN(i6[3]), .B(n25), .C(n51), .Y(r4[3]) );
  OR2X8 U73 ( .A(n46), .B(n27), .Y(n86) );
  CLKINVX40 U74 ( .A(n86), .Y(r5[1]) );
  CLKBUFX40 U75 ( .A(i5[0]), .Y(n87) );
endmodule


module sign_xor_10 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35;

  XOR2XLTH U1 ( .A(n30), .B(n24), .Y(out6) );
  XOR2XL U2 ( .A(in4), .B(n24), .Y(out4) );
  XOR2XL U3 ( .A(n32), .B(n24), .Y(out5) );
  XOR2X1 U4 ( .A(in1), .B(n24), .Y(out1) );
  CLKXOR2X4 U5 ( .A(in4), .B(n4), .Y(n3) );
  XOR2X2 U6 ( .A(n25), .B(n26), .Y(n4) );
  XNOR2X4 U8 ( .A(in1), .B(n5), .Y(n2) );
  XOR2XLTH U9 ( .A(n35), .B(n24), .Y(out2) );
  XOR2X3TH U10 ( .A(n27), .B(n28), .Y(n5) );
  XNOR2X4 U11 ( .A(n2), .B(n3), .Y(n1) );
  CLKINVX40 U7 ( .A(n1), .Y(n23) );
  CLKINVX40 U12 ( .A(n23), .Y(n24) );
  XNOR2X1 U13 ( .A(n33), .B(n24), .Y(out3) );
  DLY1X1TH U14 ( .A(in6), .Y(n25) );
  DLY1X1TH U15 ( .A(in5), .Y(n26) );
  DLY1X1TH U16 ( .A(in3), .Y(n27) );
  DLY1X1TH U17 ( .A(in2), .Y(n28) );
  INVXLTH U18 ( .A(n25), .Y(n29) );
  INVXLTH U19 ( .A(n29), .Y(n30) );
  INVXLTH U20 ( .A(n26), .Y(n31) );
  INVXLTH U21 ( .A(n31), .Y(n32) );
  INVXLTH U22 ( .A(n27), .Y(n33) );
  INVXLTH U23 ( .A(n28), .Y(n34) );
  INVXLTH U24 ( .A(n34), .Y(n35) );
endmodule


module all6_10 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100;

  sign_xor_10 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X2 U1 ( .A(n59), .B(n27), .C(n62), .Y(r4[1]) );
  NAND3X2 U3 ( .A(i6[1]), .B(n91), .C(n90), .Y(n31) );
  NOR3X1TH U4 ( .A(n60), .B(n26), .C(n64), .Y(r4[2]) );
  NOR3X1TH U5 ( .A(n30), .B(n80), .C(n75), .Y(r3[2]) );
  NOR2X2 U6 ( .A(n56), .B(n32), .Y(r1[0]) );
  NAND3X2 U7 ( .A(i6[2]), .B(n86), .C(n85), .Y(n30) );
  NOR3X1TH U8 ( .A(n64), .B(n26), .C(n68), .Y(r6[2]) );
  NOR3X4TH U9 ( .A(n63), .B(n28), .C(n67), .Y(r6[0]) );
  OR2XLTH U11 ( .A(n72), .B(n75), .Y(n52) );
  OR2X1 U13 ( .A(n76), .B(n31), .Y(n54) );
  NOR2X2 U14 ( .A(n52), .B(n30), .Y(r1[2]) );
  INVXL U15 ( .A(n89), .Y(n75) );
  INVX1 U16 ( .A(n97), .Y(n72) );
  OR2X1TH U18 ( .A(n58), .B(n67), .Y(n53) );
  NAND3X2TH U19 ( .A(n88), .B(n84), .C(n83), .Y(n25) );
  INVXLTH U20 ( .A(i6[0]), .Y(n58) );
  NOR3X4TH U21 ( .A(n58), .B(n28), .C(n63), .Y(r4[0]) );
  INVX2 U23 ( .A(n94), .Y(n74) );
  INVXLTH U24 ( .A(i3[0]), .Y(n70) );
  NAND3X4 U25 ( .A(n94), .B(i1[0]), .C(i3[0]), .Y(n28) );
  CLKINVX1TH U26 ( .A(i4[0]), .Y(n67) );
  INVX1TH U27 ( .A(n93), .Y(n78) );
  INVX1TH U28 ( .A(n91), .Y(n66) );
  CLKINVX1TH U29 ( .A(i5[0]), .Y(n63) );
  NOR3X1TH U30 ( .A(n57), .B(n25), .C(n61), .Y(r4[3]) );
  INVXLTH U31 ( .A(n87), .Y(n80) );
  INVXLTH U32 ( .A(i3[1]), .Y(n71) );
  OR2XLTH U33 ( .A(n71), .B(n76), .Y(n55) );
  OR2XLTH U34 ( .A(n70), .B(n74), .Y(n56) );
  CLKINVX1TH U35 ( .A(n90), .Y(n62) );
  NOR3X2 U36 ( .A(n59), .B(n27), .C(n66), .Y(r5[1]) );
  NOR3X1TH U37 ( .A(n61), .B(n25), .C(n65), .Y(r6[3]) );
  INVXLTH U38 ( .A(n83), .Y(n69) );
  NOR3X1TH U39 ( .A(n57), .B(n25), .C(n65), .Y(r5[3]) );
  NAND3X3TH U40 ( .A(n92), .B(n93), .C(i3[1]), .Y(n27) );
  INVXLTH U41 ( .A(i6[1]), .Y(n59) );
  NAND3X2TH U42 ( .A(i5[3]), .B(n96), .C(n95), .Y(n29) );
  INVXLTH U43 ( .A(n88), .Y(n73) );
  INVXLTH U44 ( .A(n84), .Y(n77) );
  INVX1TH U45 ( .A(n92), .Y(n76) );
  NOR3X1TH U46 ( .A(n29), .B(n73), .C(n69), .Y(r1[3]) );
  NOR3X4TH U47 ( .A(n62), .B(n27), .C(n66), .Y(r6[1]) );
  NOR3X2TH U48 ( .A(n31), .B(n78), .C(n71), .Y(r2[1]) );
  NOR3X2 U49 ( .A(n32), .B(n79), .C(n70), .Y(r2[0]) );
  INVXLTH U50 ( .A(i1[0]), .Y(n79) );
  NOR3X4TH U51 ( .A(n32), .B(n79), .C(n74), .Y(r3[0]) );
  NOR3X1TH U52 ( .A(n29), .B(n77), .C(n73), .Y(r3[3]) );
  NOR3X1TH U53 ( .A(n29), .B(n77), .C(n69), .Y(r2[3]) );
  NOR3XLTH U54 ( .A(n60), .B(n26), .C(n68), .Y(r5[2]) );
  NOR3XLTH U55 ( .A(n30), .B(n80), .C(n72), .Y(r2[2]) );
  INVXLTH U56 ( .A(i6[2]), .Y(n60) );
  INVXLTH U57 ( .A(n95), .Y(n57) );
  INVXLTH U58 ( .A(n85), .Y(n64) );
  INVXLTH U59 ( .A(i5[3]), .Y(n61) );
  INVXLTH U60 ( .A(n86), .Y(n68) );
  INVXLTH U61 ( .A(n96), .Y(n65) );
  AND3X8 U2 ( .A(n89), .B(n87), .C(n97), .Y(n81) );
  CLKINVX40 U10 ( .A(n81), .Y(n26) );
  OR2X8 U12 ( .A(n55), .B(n31), .Y(n82) );
  CLKINVX40 U17 ( .A(n82), .Y(r1[1]) );
  DLY1X1TH U22 ( .A(i3[3]), .Y(n83) );
  DLY1X1TH U62 ( .A(i1[3]), .Y(n84) );
  DLY1X1TH U63 ( .A(i5[2]), .Y(n85) );
  DLY1X1TH U64 ( .A(i4[2]), .Y(n86) );
  DLY1X1TH U65 ( .A(i1[2]), .Y(n87) );
  DLY1X1TH U66 ( .A(i2[3]), .Y(n88) );
  DLY1X1TH U67 ( .A(i2[2]), .Y(n89) );
  DLY1X1TH U68 ( .A(i5[1]), .Y(n90) );
  DLY1X1TH U69 ( .A(i4[1]), .Y(n91) );
  DLY1X1TH U70 ( .A(i2[1]), .Y(n92) );
  DLY1X1TH U71 ( .A(i1[1]), .Y(n93) );
  DLY1X1TH U72 ( .A(i2[0]), .Y(n94) );
  DLY1X1TH U73 ( .A(i6[3]), .Y(n95) );
  DLY1X1TH U74 ( .A(i4[3]), .Y(n96) );
  DLY1X1TH U75 ( .A(i3[2]), .Y(n97) );
  OR2X8 U76 ( .A(n53), .B(n28), .Y(n98) );
  CLKINVX40 U77 ( .A(n98), .Y(r5[0]) );
  OR2X8 U78 ( .A(n54), .B(n78), .Y(n99) );
  CLKINVX40 U79 ( .A(n99), .Y(r3[1]) );
  AND3X8 U80 ( .A(i5[0]), .B(i4[0]), .C(i6[0]), .Y(n100) );
  CLKINVX40 U81 ( .A(n100), .Y(n32) );
endmodule


module sign_xor_9 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n4, n5, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42;

  NAND2X5 U2 ( .A(in6), .B(n21), .Y(n22) );
  NAND2X6 U3 ( .A(n20), .B(in5), .Y(n23) );
  CLKNAND2X8 U4 ( .A(n22), .B(n23), .Y(n4) );
  INVX4 U5 ( .A(in6), .Y(n20) );
  INVX5 U6 ( .A(in5), .Y(n21) );
  INVX3 U7 ( .A(n4), .Y(n25) );
  CLKNAND2X4 U8 ( .A(in4), .B(n4), .Y(n26) );
  XOR2XL U9 ( .A(n41), .B(n37), .Y(out1) );
  CLKINVX6 U10 ( .A(in4), .Y(n24) );
  XOR2X3 U11 ( .A(in5), .B(n37), .Y(out5) );
  INVX1TH U12 ( .A(n37), .Y(n29) );
  XOR2X4TH U13 ( .A(in3), .B(in2), .Y(n5) );
  CLKNAND2X4 U14 ( .A(n26), .B(n27), .Y(n32) );
  CLKXOR2X8TH U16 ( .A(n2), .B(n32), .Y(n1) );
  XNOR2X4TH U19 ( .A(n39), .B(n5), .Y(n2) );
  NAND2X3 U20 ( .A(n24), .B(n25), .Y(n27) );
  NAND2X1TH U21 ( .A(in2), .B(n29), .Y(n30) );
  NAND2XLTH U22 ( .A(n28), .B(n37), .Y(n31) );
  INVXLTH U23 ( .A(in2), .Y(n28) );
  XNOR2X1 U1 ( .A(in4), .B(n35), .Y(out4) );
  XNOR2X1 U15 ( .A(n33), .B(n37), .Y(out6) );
  CLKINVX40 U17 ( .A(in6), .Y(n33) );
  AND2X8 U18 ( .A(n30), .B(n31), .Y(n34) );
  CLKINVX40 U24 ( .A(n34), .Y(out2) );
  CLKINVX40 U25 ( .A(n1), .Y(n35) );
  CLKINVX40 U26 ( .A(n35), .Y(n36) );
  CLKINVX40 U27 ( .A(n35), .Y(n37) );
  DLY1X1TH U28 ( .A(n42), .Y(n38) );
  DLY1X1TH U29 ( .A(in1), .Y(n39) );
  INVXLTH U30 ( .A(n39), .Y(n40) );
  INVXLTH U31 ( .A(n40), .Y(n41) );
  XNOR2X1 U32 ( .A(in3), .B(n36), .Y(n42) );
  CLKINVX40 U33 ( .A(n38), .Y(out3) );
endmodule


module all6_9 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99;

  NAND3X2 U1 ( .A(n98), .B(n97), .C(n96), .Y(n25) );
  sign_xor_9 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  INVX2 U2 ( .A(n92), .Y(n70) );
  BUFX2 U3 ( .A(n27), .Y(n54) );
  NAND3X2TH U4 ( .A(i4[2]), .B(n87), .C(n86), .Y(n30) );
  NOR2X6 U5 ( .A(n51), .B(n58), .Y(r5[0]) );
  NOR3X2 U6 ( .A(n29), .B(n78), .C(n73), .Y(r3[3]) );
  NOR3X4 U7 ( .A(n31), .B(n77), .C(n71), .Y(r3[1]) );
  INVX2 U8 ( .A(i1[1]), .Y(n77) );
  NOR3X1TH U9 ( .A(n55), .B(n25), .C(n63), .Y(r5[3]) );
  NOR3XL U10 ( .A(n30), .B(n75), .C(n74), .Y(r3[2]) );
  NOR3X1TH U11 ( .A(n57), .B(n26), .C(n64), .Y(r5[2]) );
  NOR3X1 U12 ( .A(n30), .B(n75), .C(n69), .Y(r2[2]) );
  OR2X2TH U13 ( .A(n66), .B(n28), .Y(n51) );
  INVX1TH U14 ( .A(n95), .Y(n58) );
  NAND3X4 U15 ( .A(i5[0]), .B(i4[0]), .C(n95), .Y(n32) );
  INVX2 U17 ( .A(i4[0]), .Y(n66) );
  NAND3X2TH U18 ( .A(i6[3]), .B(i4[3]), .C(n85), .Y(n29) );
  INVXLTH U19 ( .A(n97), .Y(n78) );
  NAND3X4TH U20 ( .A(i5[1]), .B(i4[1]), .C(i6[1]), .Y(n31) );
  INVX1TH U21 ( .A(n89), .Y(n71) );
  NOR3X1TH U22 ( .A(n62), .B(n26), .C(n64), .Y(r6[2]) );
  NOR3X4TH U23 ( .A(n56), .B(n54), .C(n65), .Y(r5[1]) );
  NOR3X4 U24 ( .A(n31), .B(n77), .C(n68), .Y(r2[1]) );
  INVXLTH U25 ( .A(n98), .Y(n73) );
  INVXLTH U26 ( .A(n94), .Y(n69) );
  NOR3X1TH U27 ( .A(n55), .B(n25), .C(n59), .Y(r4[3]) );
  INVXLTH U29 ( .A(n96), .Y(n67) );
  INVX1TH U30 ( .A(i5[0]), .Y(n60) );
  NAND3X2TH U31 ( .A(i1[1]), .B(n89), .C(n88), .Y(n27) );
  NAND3X3TH U32 ( .A(n93), .B(n94), .C(i1[2]), .Y(n26) );
  CLKINVX1TH U33 ( .A(n88), .Y(n68) );
  OR2XLTH U34 ( .A(n66), .B(n60), .Y(n52) );
  OR2XLTH U35 ( .A(n70), .B(n32), .Y(n53) );
  NOR3X1TH U36 ( .A(n30), .B(n74), .C(n69), .Y(r1[2]) );
  CLKINVX1TH U37 ( .A(n93), .Y(n74) );
  CLKINVX1TH U39 ( .A(n91), .Y(n72) );
  INVXLTH U40 ( .A(i4[2]), .Y(n64) );
  CLKINVX1TH U41 ( .A(i6[1]), .Y(n56) );
  CLKINVX1TH U42 ( .A(i5[1]), .Y(n61) );
  NOR3X4TH U44 ( .A(n56), .B(n54), .C(n61), .Y(r4[1]) );
  CLKINVX1TH U45 ( .A(i4[1]), .Y(n65) );
  NOR3X1TH U46 ( .A(n29), .B(n78), .C(n67), .Y(r2[3]) );
  INVX1TH U47 ( .A(n90), .Y(n76) );
  CLKINVX1TH U48 ( .A(i1[2]), .Y(n75) );
  NOR3X1TH U51 ( .A(n59), .B(n25), .C(n63), .Y(r6[3]) );
  NOR3X4TH U52 ( .A(n31), .B(n71), .C(n68), .Y(r1[1]) );
  NOR3X1TH U53 ( .A(n29), .B(n73), .C(n67), .Y(r1[3]) );
  NOR3XL U54 ( .A(n57), .B(n26), .C(n62), .Y(r4[2]) );
  INVXLTH U55 ( .A(n86), .Y(n57) );
  INVXLTH U56 ( .A(i6[3]), .Y(n55) );
  INVXLTH U57 ( .A(n87), .Y(n62) );
  INVXLTH U58 ( .A(n85), .Y(n59) );
  INVXLTH U59 ( .A(i4[3]), .Y(n63) );
  NOR3X4 U60 ( .A(n32), .B(n76), .C(n70), .Y(r2[0]) );
  OR3X8 U16 ( .A(n80), .B(n54), .C(n65), .Y(n79) );
  CLKINVX40 U28 ( .A(n79), .Y(r6[1]) );
  CLKINVX40 U38 ( .A(i5[1]), .Y(n80) );
  AND3X8 U43 ( .A(n91), .B(n90), .C(n92), .Y(n81) );
  CLKINVX40 U49 ( .A(n81), .Y(n28) );
  OR3X8 U50 ( .A(n32), .B(n76), .C(n72), .Y(n82) );
  CLKINVX40 U61 ( .A(n82), .Y(r3[0]) );
  OR3X8 U62 ( .A(n58), .B(n28), .C(n60), .Y(n83) );
  CLKINVX40 U63 ( .A(n83), .Y(r4[0]) );
  OR2X8 U64 ( .A(n53), .B(n72), .Y(n84) );
  CLKINVX40 U65 ( .A(n84), .Y(r1[0]) );
  DLY1X1TH U66 ( .A(i5[3]), .Y(n85) );
  DLY1X1TH U67 ( .A(i6[2]), .Y(n86) );
  DLY1X1TH U68 ( .A(i5[2]), .Y(n87) );
  DLY1X1TH U69 ( .A(i3[1]), .Y(n88) );
  DLY1X1TH U70 ( .A(i2[1]), .Y(n89) );
  DLY1X1TH U71 ( .A(i1[0]), .Y(n90) );
  DLY1X1TH U72 ( .A(i2[0]), .Y(n91) );
  DLY1X1TH U73 ( .A(i3[0]), .Y(n92) );
  DLY1X1TH U74 ( .A(i2[2]), .Y(n93) );
  DLY1X1TH U75 ( .A(i3[2]), .Y(n94) );
  DLY1X1TH U76 ( .A(i6[0]), .Y(n95) );
  DLY1X1TH U77 ( .A(i3[3]), .Y(n96) );
  DLY1X1TH U78 ( .A(i1[3]), .Y(n97) );
  DLY1X1TH U79 ( .A(i2[3]), .Y(n98) );
  OR2X8 U80 ( .A(n52), .B(n28), .Y(n99) );
  CLKINVX40 U81 ( .A(n99), .Y(r6[0]) );
endmodule


module sign_xor_8 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n27, n28, n29, n30, n31, n32, n33, n34, n35;

  XOR2X1 U1 ( .A(in3), .B(in2), .Y(n5) );
  XOR2X1 U2 ( .A(in4), .B(n31), .Y(out4) );
  BUFX16 U3 ( .A(n1), .Y(n31) );
  XOR2X1 U4 ( .A(in6), .B(n31), .Y(out6) );
  CLKNAND2X4 U5 ( .A(in1), .B(n28), .Y(n29) );
  CLKNAND2X2 U6 ( .A(n27), .B(n31), .Y(n30) );
  NAND2X8 U7 ( .A(n29), .B(n30), .Y(out1) );
  INVX1TH U8 ( .A(in1), .Y(n27) );
  INVX1 U9 ( .A(n31), .Y(n28) );
  XOR2XLTH U10 ( .A(in2), .B(n31), .Y(out2) );
  CLKNAND2X4 U11 ( .A(n34), .B(n35), .Y(out5) );
  XOR2X1 U12 ( .A(in6), .B(in5), .Y(n4) );
  NAND2XLTH U13 ( .A(n32), .B(n31), .Y(n35) );
  XOR2X1 U14 ( .A(in3), .B(n31), .Y(out3) );
  XNOR2X4 U15 ( .A(in1), .B(n5), .Y(n2) );
  INVX2TH U16 ( .A(n31), .Y(n33) );
  XOR2X8 U17 ( .A(n4), .B(in4), .Y(n3) );
  CLKNAND2X2 U18 ( .A(in5), .B(n33), .Y(n34) );
  INVXLTH U19 ( .A(in5), .Y(n32) );
  XNOR2X4 U20 ( .A(n2), .B(n3), .Y(n1) );
endmodule


module all6_8 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92;

  NOR3X1 U50 ( .A(n30), .B(n69), .C(n61), .Y(r2[2]) );
  sign_xor_8 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X2 U2 ( .A(n31), .B(n66), .C(n60), .Y(r2[1]) );
  NOR3XL U3 ( .A(n32), .B(n67), .C(n59), .Y(r2[0]) );
  NOR3X1 U5 ( .A(n31), .B(n66), .C(n62), .Y(r3[1]) );
  INVX1TH U7 ( .A(i4[0]), .Y(n56) );
  NAND3X4TH U8 ( .A(n81), .B(n82), .C(i1[2]), .Y(n26) );
  NOR3X1TH U9 ( .A(n49), .B(n26), .C(n51), .Y(r4[2]) );
  NOR3X4 U10 ( .A(n53), .B(n27), .C(n55), .Y(r6[1]) );
  NAND3X2 U11 ( .A(i4[2]), .B(n79), .C(n77), .Y(n30) );
  NOR3X2 U12 ( .A(n31), .B(n62), .C(n60), .Y(r1[1]) );
  INVXLTH U14 ( .A(i5[3]), .Y(n50) );
  NOR3X1TH U15 ( .A(n47), .B(n25), .C(n86), .Y(r4[3]) );
  NOR3X1TH U16 ( .A(n49), .B(n26), .C(n57), .Y(r5[2]) );
  INVXLTH U17 ( .A(i1[3]), .Y(n68) );
  INVXLTH U19 ( .A(i4[2]), .Y(n57) );
  CLKINVX1TH U20 ( .A(i5[1]), .Y(n53) );
  INVXLTH U22 ( .A(i3[0]), .Y(n59) );
  NOR3X1TH U23 ( .A(n65), .B(n69), .C(n30), .Y(r3[2]) );
  NOR3X1TH U24 ( .A(n32), .B(n88), .C(n59), .Y(r1[0]) );
  NOR2X6TH U25 ( .A(n45), .B(n48), .Y(r5[0]) );
  INVXLTH U26 ( .A(n76), .Y(n58) );
  INVX1TH U27 ( .A(i6[0]), .Y(n48) );
  INVX2TH U28 ( .A(n85), .Y(n52) );
  NOR3X1TH U29 ( .A(n29), .B(n64), .C(n58), .Y(r1[3]) );
  INVXLTH U30 ( .A(n75), .Y(n54) );
  INVXLTH U31 ( .A(n77), .Y(n49) );
  NAND3X4TH U33 ( .A(n85), .B(i4[0]), .C(i6[0]), .Y(n32) );
  OR2XLTH U34 ( .A(n56), .B(n28), .Y(n45) );
  INVX1TH U35 ( .A(n84), .Y(n55) );
  NOR3X1TH U36 ( .A(n29), .B(n68), .C(n58), .Y(r2[3]) );
  NOR3X4 U37 ( .A(n52), .B(n28), .C(n56), .Y(r6[0]) );
  INVXLTH U38 ( .A(n80), .Y(n64) );
  INVXLTH U39 ( .A(n74), .Y(n47) );
  INVXLTH U40 ( .A(n79), .Y(n51) );
  INVX1TH U41 ( .A(n83), .Y(n46) );
  NOR3X1TH U42 ( .A(n29), .B(n68), .C(n64), .Y(r3[3]) );
  INVXLTH U43 ( .A(i1[2]), .Y(n69) );
  CLKINVX1TH U44 ( .A(i1[1]), .Y(n66) );
  INVXLTH U45 ( .A(n82), .Y(n61) );
  INVXLTH U46 ( .A(i2[0]), .Y(n63) );
  NOR3X1TH U47 ( .A(n47), .B(n25), .C(n54), .Y(r5[3]) );
  NOR3X1TH U48 ( .A(n51), .B(n26), .C(n57), .Y(r6[2]) );
  NOR3XLTH U52 ( .A(n30), .B(n65), .C(n61), .Y(r1[2]) );
  NAND3X4 U53 ( .A(i2[0]), .B(i1[0]), .C(i3[0]), .Y(n28) );
  INVXLTH U54 ( .A(i2[1]), .Y(n62) );
  INVXLTH U55 ( .A(n81), .Y(n65) );
  INVXLTH U56 ( .A(n78), .Y(n60) );
  CLKINVX1TH U57 ( .A(i1[0]), .Y(n67) );
  AND3X8 U1 ( .A(i5[3]), .B(n75), .C(n74), .Y(n70) );
  CLKINVX40 U4 ( .A(n70), .Y(n29) );
  AND3X8 U6 ( .A(i1[3]), .B(n80), .C(n76), .Y(n71) );
  CLKINVX40 U13 ( .A(n71), .Y(n25) );
  NOR3BX4 U18 ( .AN(i6[0]), .B(n28), .C(n52), .Y(r4[0]) );
  AND3X8 U21 ( .A(i2[1]), .B(i1[1]), .C(n78), .Y(n72) );
  CLKINVX40 U32 ( .A(n72), .Y(n27) );
  OR3X8 U49 ( .A(n46), .B(n27), .C(n55), .Y(n73) );
  CLKINVX40 U51 ( .A(n73), .Y(r5[1]) );
  DLY1X1TH U58 ( .A(i6[3]), .Y(n74) );
  DLY1X1TH U59 ( .A(i4[3]), .Y(n75) );
  DLY1X1TH U60 ( .A(i3[3]), .Y(n76) );
  DLY1X1TH U61 ( .A(i6[2]), .Y(n77) );
  DLY1X1TH U62 ( .A(i3[1]), .Y(n78) );
  DLY1X1TH U63 ( .A(i5[2]), .Y(n79) );
  DLY1X1TH U64 ( .A(i2[3]), .Y(n80) );
  DLY1X1TH U65 ( .A(i2[2]), .Y(n81) );
  DLY1X1TH U66 ( .A(i3[2]), .Y(n82) );
  DLY1X1TH U67 ( .A(i6[1]), .Y(n83) );
  DLY1X1TH U68 ( .A(i4[1]), .Y(n84) );
  DLY1X1TH U69 ( .A(i5[0]), .Y(n85) );
  INVXLTH U70 ( .A(i5[3]), .Y(n86) );
  DLY1X1TH U71 ( .A(n54), .Y(n87) );
  INVXLTH U72 ( .A(i2[0]), .Y(n88) );
  OR3X8 U73 ( .A(n32), .B(n67), .C(n63), .Y(n89) );
  CLKINVX40 U74 ( .A(n89), .Y(r3[0]) );
  OR3X8 U75 ( .A(n46), .B(n27), .C(n53), .Y(n90) );
  CLKINVX40 U76 ( .A(n90), .Y(r4[1]) );
  AND3X8 U77 ( .A(i5[1]), .B(n84), .C(n83), .Y(n91) );
  CLKINVX40 U78 ( .A(n91), .Y(n31) );
  OR3X8 U79 ( .A(n50), .B(n25), .C(n87), .Y(n92) );
  CLKINVX40 U80 ( .A(n92), .Y(r6[3]) );
endmodule


module sign_xor_7 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n3, n4, n5, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38;

  CLKNAND2X4 U1 ( .A(n25), .B(n26), .Y(out3) );
  NAND2X4 U2 ( .A(n29), .B(n30), .Y(out2) );
  XOR2X1 U3 ( .A(n38), .B(n1), .Y(out1) );
  NAND2XLTH U4 ( .A(in3), .B(n28), .Y(n25) );
  NAND2XLTH U5 ( .A(n24), .B(n1), .Y(n26) );
  INVX2TH U6 ( .A(n1), .Y(n28) );
  XOR2X4 U7 ( .A(n34), .B(n5), .Y(n31) );
  XOR2X3 U8 ( .A(n33), .B(n4), .Y(n3) );
  INVXLTH U9 ( .A(in3), .Y(n24) );
  XOR2X8 U10 ( .A(n31), .B(n3), .Y(n1) );
  XOR2X3TH U11 ( .A(in3), .B(in2), .Y(n5) );
  XOR2XLTH U12 ( .A(in5), .B(n1), .Y(out5) );
  XOR2X1TH U13 ( .A(n36), .B(n1), .Y(out4) );
  NAND2XLTH U15 ( .A(n27), .B(n1), .Y(n30) );
  INVXLTH U16 ( .A(in2), .Y(n27) );
  XOR2X1TH U17 ( .A(in6), .B(n1), .Y(out6) );
  XOR2X2 U18 ( .A(in6), .B(in5), .Y(n4) );
  AND2X8 U14 ( .A(in2), .B(n28), .Y(n32) );
  CLKINVX40 U19 ( .A(n32), .Y(n29) );
  DLY1X1TH U20 ( .A(in4), .Y(n33) );
  DLY1X1TH U21 ( .A(in1), .Y(n34) );
  INVXLTH U22 ( .A(n33), .Y(n35) );
  INVXLTH U23 ( .A(n35), .Y(n36) );
  INVXLTH U24 ( .A(n34), .Y(n37) );
  INVXLTH U25 ( .A(n37), .Y(n38) );
endmodule


module all6_7 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77;

  NOR3X1 U38 ( .A(n42), .B(n26), .C(n51), .Y(r5[2]) );
  sign_xor_7 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X1 U1 ( .A(n30), .B(n58), .C(n54), .Y(r1[2]) );
  NOR2X4 U2 ( .A(n44), .B(n28), .Y(n35) );
  NOR2X4 U3 ( .A(n36), .B(n49), .Y(r5[0]) );
  INVX2 U4 ( .A(n35), .Y(n36) );
  NAND3X4 U5 ( .A(n75), .B(i1[0]), .C(i2[0]), .Y(n28) );
  NOR3X1 U7 ( .A(n32), .B(n64), .C(n60), .Y(r3[0]) );
  OR2XLTH U8 ( .A(n55), .B(n31), .Y(n37) );
  INVX2 U9 ( .A(i6[0]), .Y(n44) );
  NOR2X4 U10 ( .A(n37), .B(n59), .Y(r1[1]) );
  INVX1 U11 ( .A(n74), .Y(n59) );
  CLKINVX2 U12 ( .A(i3[1]), .Y(n55) );
  NAND3X4 U14 ( .A(i2[2]), .B(i1[2]), .C(i3[2]), .Y(n26) );
  INVXLTH U15 ( .A(i2[0]), .Y(n60) );
  NOR2X6 U16 ( .A(n31), .B(n63), .Y(n38) );
  NOR2X4 U17 ( .A(n39), .B(n55), .Y(r2[1]) );
  INVX6TH U18 ( .A(n38), .Y(n39) );
  CLKINVX1 U19 ( .A(i1[1]), .Y(n63) );
  NAND3X3TH U20 ( .A(n70), .B(i1[1]), .C(i3[1]), .Y(n27) );
  INVXLTH U21 ( .A(i3[2]), .Y(n54) );
  NOR3X4TH U22 ( .A(n29), .B(n57), .C(n56), .Y(r1[3]) );
  NOR3X1TH U23 ( .A(n42), .B(n26), .C(n46), .Y(r4[2]) );
  NOR3X1TH U24 ( .A(n30), .B(n62), .C(n58), .Y(r3[2]) );
  NOR3XL U25 ( .A(n30), .B(n62), .C(n54), .Y(r2[2]) );
  CLKINVX1TH U26 ( .A(i1[0]), .Y(n64) );
  INVXLTH U28 ( .A(i5[2]), .Y(n46) );
  NAND3X2TH U29 ( .A(i5[2]), .B(i4[2]), .C(i6[2]), .Y(n30) );
  NOR2X4TH U30 ( .A(n40), .B(n53), .Y(r1[0]) );
  OR2XLTH U31 ( .A(n60), .B(n32), .Y(n40) );
  NOR3X2 U32 ( .A(n43), .B(n27), .C(n47), .Y(r4[1]) );
  CLKINVX1TH U33 ( .A(n73), .Y(n52) );
  INVXLTH U34 ( .A(i6[2]), .Y(n42) );
  NOR3X4TH U35 ( .A(n47), .B(n27), .C(n52), .Y(r6[1]) );
  INVXLTH U36 ( .A(n68), .Y(n50) );
  INVXLTH U37 ( .A(n69), .Y(n61) );
  INVXLTH U39 ( .A(n67), .Y(n56) );
  INVXLTH U40 ( .A(i2[3]), .Y(n57) );
  NAND3X2TH U41 ( .A(i2[3]), .B(n69), .C(n67), .Y(n25) );
  INVXLTH U42 ( .A(i6[3]), .Y(n41) );
  INVXLTH U43 ( .A(i5[3]), .Y(n45) );
  NOR3X1TH U44 ( .A(n45), .B(n25), .C(n50), .Y(r6[3]) );
  INVXLTH U45 ( .A(i4[2]), .Y(n51) );
  NOR3X1TH U46 ( .A(n41), .B(n25), .C(n50), .Y(r5[3]) );
  INVXLTH U47 ( .A(i6[1]), .Y(n43) );
  NOR3X1TH U48 ( .A(n29), .B(n61), .C(n57), .Y(r3[3]) );
  NOR3X1TH U49 ( .A(n29), .B(n61), .C(n56), .Y(r2[3]) );
  NOR3X1TH U50 ( .A(n41), .B(n25), .C(n45), .Y(r4[3]) );
  NOR3XLTH U51 ( .A(n46), .B(n26), .C(n51), .Y(r6[2]) );
  NOR3X4TH U52 ( .A(n43), .B(n27), .C(n52), .Y(r5[1]) );
  NOR3X4 U53 ( .A(n32), .B(n64), .C(n53), .Y(r2[0]) );
  CLKINVX1TH U54 ( .A(n71), .Y(n48) );
  INVX2 U56 ( .A(n75), .Y(n53) );
  CLKINVX1TH U57 ( .A(n72), .Y(n49) );
  NAND3X4 U58 ( .A(n71), .B(n72), .C(n77), .Y(n32) );
  INVXLTH U59 ( .A(i5[1]), .Y(n47) );
  NOR3X2 U60 ( .A(n31), .B(n63), .C(n59), .Y(r3[1]) );
  INVXLTH U61 ( .A(i1[2]), .Y(n62) );
  INVXLTH U62 ( .A(i2[2]), .Y(n58) );
  AND3X8 U6 ( .A(i5[3]), .B(n68), .C(i6[3]), .Y(n65) );
  CLKINVX40 U13 ( .A(n65), .Y(n29) );
  NOR3X8 U27 ( .A(n44), .B(n28), .C(n48), .Y(r4[0]) );
  AND3X8 U55 ( .A(i5[1]), .B(n73), .C(i6[1]), .Y(n66) );
  CLKINVX40 U63 ( .A(n66), .Y(n31) );
  DLY1X1TH U64 ( .A(i3[3]), .Y(n67) );
  DLY1X1TH U65 ( .A(i4[3]), .Y(n68) );
  DLY1X1TH U66 ( .A(i1[3]), .Y(n69) );
  DLY1X1TH U67 ( .A(i2[1]), .Y(n70) );
  DLY1X1TH U68 ( .A(i5[0]), .Y(n71) );
  DLY1X1TH U69 ( .A(i4[0]), .Y(n72) );
  DLY1X1TH U70 ( .A(i4[1]), .Y(n73) );
  DLY1X1TH U71 ( .A(n70), .Y(n74) );
  DLY1X1TH U72 ( .A(i3[0]), .Y(n75) );
  OR3X8 U73 ( .A(n48), .B(n28), .C(n49), .Y(n76) );
  CLKINVX40 U74 ( .A(n76), .Y(r6[0]) );
  CLKINVX40 U75 ( .A(n44), .Y(n77) );
endmodule


module sign_xor_6 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33;

  XOR2X1 U1 ( .A(in6), .B(in5), .Y(n4) );
  CLKXOR2X4 U2 ( .A(n4), .B(n31), .Y(n3) );
  XNOR2X4 U3 ( .A(in1), .B(n5), .Y(n2) );
  NAND2X1 U4 ( .A(in3), .B(n23), .Y(n24) );
  NAND2XL U5 ( .A(n22), .B(n26), .Y(n25) );
  CLKNAND2X4 U6 ( .A(n24), .B(n25), .Y(out3) );
  CLKINVX2TH U7 ( .A(in3), .Y(n22) );
  INVX4 U8 ( .A(n26), .Y(n23) );
  BUFX20 U9 ( .A(n1), .Y(n26) );
  CLKNAND2X4 U10 ( .A(n29), .B(n30), .Y(out1) );
  XOR2X2TH U11 ( .A(in3), .B(in2), .Y(n5) );
  NAND2XLTH U12 ( .A(in1), .B(n28), .Y(n29) );
  XOR2XL U13 ( .A(n33), .B(n26), .Y(out4) );
  INVXLTH U14 ( .A(n26), .Y(n28) );
  XOR2XLTH U15 ( .A(in5), .B(n26), .Y(out5) );
  NAND2X2 U16 ( .A(n27), .B(n26), .Y(n30) );
  INVXLTH U17 ( .A(in1), .Y(n27) );
  XOR2X1TH U18 ( .A(in2), .B(n26), .Y(out2) );
  XOR2X1TH U19 ( .A(in6), .B(n26), .Y(out6) );
  XNOR2X4 U20 ( .A(n2), .B(n3), .Y(n1) );
  DLY1X1TH U21 ( .A(in4), .Y(n31) );
  INVXLTH U22 ( .A(n31), .Y(n32) );
  INVXLTH U23 ( .A(n32), .Y(n33) );
endmodule


module all6_6 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98;

  NAND3X2 U6 ( .A(n97), .B(n96), .C(n95), .Y(n30) );
  sign_xor_6 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X2 U1 ( .A(n58), .B(n28), .C(n67), .Y(r5[0]) );
  INVXL U2 ( .A(i1[0]), .Y(n78) );
  NOR2X4 U4 ( .A(n55), .B(n75), .Y(r1[0]) );
  OR2XLTH U5 ( .A(n76), .B(n92), .Y(n53) );
  NOR3X1 U7 ( .A(n30), .B(n77), .C(n71), .Y(r2[2]) );
  INVX2 U8 ( .A(n90), .Y(n71) );
  NOR3X4 U9 ( .A(n60), .B(n27), .C(n65), .Y(r6[1]) );
  NAND3X2 U10 ( .A(i2[1]), .B(i1[1]), .C(i3[1]), .Y(n27) );
  NOR2X4 U11 ( .A(n53), .B(n29), .Y(r3[3]) );
  NOR2X2 U12 ( .A(n32), .B(n70), .Y(n54) );
  CLKINVX2 U13 ( .A(n54), .Y(n55) );
  INVX2 U14 ( .A(i2[0]), .Y(n75) );
  INVX2 U15 ( .A(i3[0]), .Y(n70) );
  NOR3X2 U16 ( .A(n30), .B(n73), .C(n71), .Y(r1[2]) );
  NOR3X4 U18 ( .A(n57), .B(n27), .C(n60), .Y(r4[1]) );
  NOR3XL U19 ( .A(n32), .B(n78), .C(n70), .Y(r2[0]) );
  NOR3X4 U20 ( .A(n30), .B(n77), .C(n73), .Y(r3[2]) );
  INVXLTH U21 ( .A(n96), .Y(n66) );
  INVX1TH U22 ( .A(i4[1]), .Y(n65) );
  NAND3X4TH U23 ( .A(n89), .B(n90), .C(i1[2]), .Y(n26) );
  CLKINVX1TH U24 ( .A(n87), .Y(n57) );
  CLKINVX1TH U25 ( .A(n88), .Y(n60) );
  NOR3X2TH U26 ( .A(n56), .B(n25), .C(n61), .Y(r4[3]) );
  NOR3X4 U27 ( .A(n58), .B(n28), .C(n63), .Y(r4[0]) );
  NOR3X1 U28 ( .A(n81), .B(n26), .C(n66), .Y(r5[2]) );
  NOR3X4 U29 ( .A(n63), .B(n28), .C(n67), .Y(r6[0]) );
  NOR3X4TH U30 ( .A(n56), .B(n25), .C(n64), .Y(r5[3]) );
  NOR3X4 U31 ( .A(n32), .B(n78), .C(n75), .Y(r3[0]) );
  INVXLTH U33 ( .A(i3[3]), .Y(n68) );
  INVXLTH U34 ( .A(i2[3]), .Y(n72) );
  INVXLTH U35 ( .A(n86), .Y(n61) );
  NAND3X2TH U36 ( .A(i3[3]), .B(n94), .C(i2[3]), .Y(n25) );
  INVXLTH U37 ( .A(n84), .Y(n56) );
  NOR3X4TH U38 ( .A(n57), .B(n27), .C(n65), .Y(r5[1]) );
  CLKINVX1TH U39 ( .A(i2[1]), .Y(n74) );
  NOR3X4 U40 ( .A(n81), .B(n26), .C(n80), .Y(r4[2]) );
  NOR3X4TH U41 ( .A(n31), .B(n79), .C(n74), .Y(r3[1]) );
  INVXLTH U42 ( .A(n85), .Y(n64) );
  INVXLTH U43 ( .A(n94), .Y(n76) );
  INVX1TH U44 ( .A(i5[0]), .Y(n63) );
  NOR3X1TH U45 ( .A(n61), .B(n25), .C(n64), .Y(r6[3]) );
  INVXLTH U46 ( .A(n95), .Y(n59) );
  NOR3X1TH U47 ( .A(n29), .B(n76), .C(n68), .Y(r2[3]) );
  NAND3X3TH U48 ( .A(i2[0]), .B(i1[0]), .C(i3[0]), .Y(n28) );
  INVX1TH U49 ( .A(n91), .Y(n67) );
  INVXLTH U50 ( .A(i6[0]), .Y(n58) );
  NOR3X4TH U51 ( .A(n31), .B(n74), .C(n69), .Y(r1[1]) );
  NOR3X2 U52 ( .A(n31), .B(n79), .C(n69), .Y(r2[1]) );
  NAND3X4 U53 ( .A(n91), .B(i5[0]), .C(i6[0]), .Y(n32) );
  INVXLTH U54 ( .A(i1[1]), .Y(n79) );
  NOR3XLTH U55 ( .A(n80), .B(n26), .C(n66), .Y(r6[2]) );
  INVXLTH U56 ( .A(i1[2]), .Y(n77) );
  INVXLTH U57 ( .A(n97), .Y(n62) );
  INVXLTH U58 ( .A(n89), .Y(n73) );
  INVXLTH U59 ( .A(i3[1]), .Y(n69) );
  CLKBUFX40 U3 ( .A(n62), .Y(n80) );
  CLKBUFX40 U17 ( .A(n59), .Y(n81) );
  AND3X8 U32 ( .A(n86), .B(n85), .C(n84), .Y(n82) );
  CLKINVX40 U60 ( .A(n82), .Y(n29) );
  AND3X8 U61 ( .A(i4[1]), .B(n88), .C(n87), .Y(n83) );
  CLKINVX40 U62 ( .A(n83), .Y(n31) );
  DLY1X1TH U63 ( .A(i6[3]), .Y(n84) );
  DLY1X1TH U64 ( .A(i4[3]), .Y(n85) );
  DLY1X1TH U65 ( .A(i5[3]), .Y(n86) );
  DLY1X1TH U66 ( .A(i6[1]), .Y(n87) );
  DLY1X1TH U67 ( .A(i5[1]), .Y(n88) );
  DLY1X1TH U68 ( .A(i2[2]), .Y(n89) );
  DLY1X1TH U69 ( .A(i3[2]), .Y(n90) );
  DLY1X1TH U70 ( .A(i4[0]), .Y(n91) );
  DLY1X1TH U71 ( .A(n72), .Y(n92) );
  DLY1X1TH U72 ( .A(n68), .Y(n93) );
  DLY1X1TH U73 ( .A(i1[3]), .Y(n94) );
  DLY1X1TH U74 ( .A(i6[2]), .Y(n95) );
  DLY1X1TH U75 ( .A(i4[2]), .Y(n96) );
  DLY1X1TH U76 ( .A(i5[2]), .Y(n97) );
  OR3X8 U77 ( .A(n29), .B(n92), .C(n93), .Y(n98) );
  CLKINVX40 U78 ( .A(n98), .Y(r1[3]) );
endmodule


module sign_xor_5 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37;

  NAND2X2 U1 ( .A(in3), .B(n30), .Y(n31) );
  NAND2X6 U2 ( .A(n27), .B(n28), .Y(n1) );
  NAND2X4 U3 ( .A(n31), .B(n32), .Y(out3) );
  XOR2X4 U4 ( .A(n37), .B(n1), .Y(out1) );
  XOR2X2 U5 ( .A(in6), .B(n1), .Y(out6) );
  XOR2X3 U6 ( .A(in3), .B(in2), .Y(n5) );
  XOR2X1 U7 ( .A(in2), .B(n1), .Y(out2) );
  INVX2 U8 ( .A(n3), .Y(n26) );
  XOR2X2 U9 ( .A(n33), .B(n4), .Y(n3) );
  INVX2TH U10 ( .A(n2), .Y(n25) );
  NAND2X2TH U11 ( .A(n2), .B(n3), .Y(n27) );
  XOR2X4 U12 ( .A(in6), .B(in5), .Y(n4) );
  XNOR2X4 U13 ( .A(in1), .B(n5), .Y(n2) );
  XOR2XL U14 ( .A(n35), .B(n1), .Y(out4) );
  XOR2XL U15 ( .A(in5), .B(n1), .Y(out5) );
  INVXLTH U16 ( .A(n1), .Y(n30) );
  NAND2X4TH U17 ( .A(n25), .B(n26), .Y(n28) );
  NAND2X1 U18 ( .A(n29), .B(n1), .Y(n32) );
  INVXLTH U19 ( .A(in3), .Y(n29) );
  DLY1X1TH U20 ( .A(in4), .Y(n33) );
  INVXLTH U21 ( .A(n33), .Y(n34) );
  INVXLTH U22 ( .A(n34), .Y(n35) );
  INVXLTH U23 ( .A(in1), .Y(n36) );
  INVXLTH U24 ( .A(n36), .Y(n37) );
endmodule


module all6_5 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82;

  NOR3X1 U34 ( .A(n49), .B(n26), .C(n54), .Y(r6[2]) );
  sign_xor_5 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X1 U1 ( .A(n30), .B(n67), .C(n59), .Y(r2[2]) );
  NOR3X1TH U2 ( .A(n46), .B(n26), .C(n54), .Y(r5[2]) );
  NOR3X4TH U3 ( .A(n47), .B(n28), .C(n55), .Y(r5[0]) );
  NAND3X2 U4 ( .A(i5[2]), .B(n75), .C(i6[2]), .Y(n30) );
  NAND3X3TH U5 ( .A(n78), .B(n79), .C(i6[3]), .Y(n29) );
  NOR3X1TH U7 ( .A(n45), .B(n25), .C(n53), .Y(r5[3]) );
  INVXLTH U8 ( .A(n78), .Y(n51) );
  NAND3X2TH U9 ( .A(i2[3]), .B(i1[3]), .C(i3[3]), .Y(n25) );
  NAND3X3TH U10 ( .A(i2[1]), .B(i1[1]), .C(i3[1]), .Y(n27) );
  INVXLTH U11 ( .A(i3[2]), .Y(n59) );
  CLKINVX1TH U12 ( .A(i2[1]), .Y(n62) );
  NOR2X4TH U13 ( .A(n43), .B(n28), .Y(r6[0]) );
  NAND3X3TH U15 ( .A(i5[0]), .B(i4[0]), .C(i6[0]), .Y(n32) );
  OR2XLTH U16 ( .A(n52), .B(n55), .Y(n43) );
  OR2XLTH U17 ( .A(n68), .B(n31), .Y(n44) );
  INVX1TH U19 ( .A(n76), .Y(n65) );
  NOR2X3 U21 ( .A(n44), .B(n62), .Y(r3[1]) );
  NAND3X4 U22 ( .A(i5[1]), .B(n81), .C(i6[1]), .Y(n31) );
  INVX1 U23 ( .A(i5[0]), .Y(n52) );
  INVX1 U25 ( .A(i4[0]), .Y(n55) );
  NOR3X1TH U26 ( .A(n29), .B(n66), .C(n57), .Y(r2[3]) );
  INVXLTH U27 ( .A(i1[3]), .Y(n66) );
  INVXLTH U28 ( .A(i2[3]), .Y(n64) );
  INVXLTH U29 ( .A(n79), .Y(n53) );
  NOR3X1TH U30 ( .A(n29), .B(n66), .C(n64), .Y(r3[3]) );
  NOR3X4TH U31 ( .A(n31), .B(n62), .C(n58), .Y(r1[1]) );
  NOR3X2 U32 ( .A(n48), .B(n27), .C(n50), .Y(r4[1]) );
  NOR3X4 U33 ( .A(n30), .B(n67), .C(n61), .Y(r3[2]) );
  NOR3X1TH U35 ( .A(n51), .B(n25), .C(n53), .Y(r6[3]) );
  INVXLTH U36 ( .A(i3[3]), .Y(n57) );
  INVXLTH U37 ( .A(n81), .Y(n56) );
  INVXLTH U38 ( .A(i6[2]), .Y(n46) );
  INVXLTH U40 ( .A(i5[2]), .Y(n49) );
  INVXLTH U41 ( .A(i5[1]), .Y(n50) );
  INVXLTH U42 ( .A(i6[3]), .Y(n45) );
  INVXLTH U43 ( .A(i3[1]), .Y(n58) );
  NOR3X1TH U44 ( .A(n29), .B(n64), .C(n57), .Y(r1[3]) );
  INVX2TH U45 ( .A(n77), .Y(n63) );
  NOR3X4TH U46 ( .A(n50), .B(n27), .C(n56), .Y(r6[1]) );
  NOR3XLTH U47 ( .A(n46), .B(n26), .C(n49), .Y(r4[2]) );
  NOR3X1TH U48 ( .A(n45), .B(n25), .C(n51), .Y(r4[3]) );
  NOR3X4TH U49 ( .A(n32), .B(n65), .C(n63), .Y(r3[0]) );
  NOR3X2 U50 ( .A(n48), .B(n27), .C(n56), .Y(r5[1]) );
  NOR3X2 U51 ( .A(n31), .B(n68), .C(n58), .Y(r2[1]) );
  INVXLTH U52 ( .A(n74), .Y(n60) );
  CLKINVX1TH U53 ( .A(i6[0]), .Y(n47) );
  INVXLTH U54 ( .A(i6[1]), .Y(n48) );
  INVXLTH U55 ( .A(i1[2]), .Y(n67) );
  INVXLTH U56 ( .A(i2[2]), .Y(n61) );
  INVXLTH U57 ( .A(i1[1]), .Y(n68) );
  INVXLTH U58 ( .A(n75), .Y(n54) );
  NOR3BX4 U6 ( .AN(n69), .B(n65), .C(n73), .Y(r2[0]) );
  CLKINVX40 U14 ( .A(n32), .Y(n69) );
  NAND3BX4 U18 ( .AN(n30), .B(i2[2]), .C(i3[2]), .Y(n70) );
  CLKINVX40 U20 ( .A(n70), .Y(r1[2]) );
  AND3X8 U24 ( .A(i2[2]), .B(i1[2]), .C(i3[2]), .Y(n71) );
  CLKINVX40 U39 ( .A(n71), .Y(n26) );
  AND3X8 U59 ( .A(n77), .B(n76), .C(n74), .Y(n72) );
  CLKINVX40 U60 ( .A(n72), .Y(n28) );
  INVXLTH U61 ( .A(n74), .Y(n73) );
  DLY1X1TH U62 ( .A(i3[0]), .Y(n74) );
  DLY1X1TH U63 ( .A(i4[2]), .Y(n75) );
  DLY1X1TH U64 ( .A(i1[0]), .Y(n76) );
  DLY1X1TH U65 ( .A(i2[0]), .Y(n77) );
  DLY1X1TH U66 ( .A(i5[3]), .Y(n78) );
  DLY1X1TH U67 ( .A(i4[3]), .Y(n79) );
  OR3X8 U68 ( .A(n60), .B(n63), .C(n32), .Y(n80) );
  CLKINVX40 U69 ( .A(n80), .Y(r1[0]) );
  CLKBUFX40 U70 ( .A(i4[1]), .Y(n81) );
  OR3X8 U71 ( .A(n47), .B(n28), .C(n52), .Y(n82) );
  CLKINVX40 U72 ( .A(n82), .Y(r4[0]) );
endmodule


module sign_xor_4 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n23, n24, n25, n26, n27, n28, n29, n30;

  CLKXOR2X2 U1 ( .A(n30), .B(n1), .Y(out1) );
  XOR2XL U2 ( .A(in6), .B(n1), .Y(out6) );
  XOR2XL U3 ( .A(in3), .B(n1), .Y(out3) );
  XOR2X3 U4 ( .A(in4), .B(n4), .Y(n3) );
  CLKXOR2X4 U5 ( .A(in6), .B(in5), .Y(n4) );
  INVX4 U6 ( .A(n3), .Y(n24) );
  CLKNAND2X8 U7 ( .A(n23), .B(n24), .Y(n26) );
  INVX4TH U8 ( .A(n2), .Y(n23) );
  XOR2XL U9 ( .A(in2), .B(n1), .Y(out2) );
  NAND2X8 U10 ( .A(n25), .B(n26), .Y(n1) );
  CLKXOR2X1TH U11 ( .A(in5), .B(n1), .Y(out5) );
  NAND2X4 U12 ( .A(n2), .B(n3), .Y(n25) );
  CLKXOR2X2TH U13 ( .A(in3), .B(in2), .Y(n5) );
  XOR2X1TH U14 ( .A(n28), .B(n1), .Y(out4) );
  XNOR2X4 U15 ( .A(in1), .B(n5), .Y(n2) );
  INVXLTH U16 ( .A(in4), .Y(n27) );
  INVXLTH U17 ( .A(n27), .Y(n28) );
  INVXLTH U18 ( .A(in1), .Y(n29) );
  INVXLTH U19 ( .A(n29), .Y(n30) );
endmodule


module all6_4 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100;

  NOR3X1 U34 ( .A(n60), .B(n26), .C(n67), .Y(r6[2]) );
  sign_xor_4 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NAND3X2 U1 ( .A(i2[1]), .B(i1[1]), .C(i3[1]), .Y(n27) );
  NAND3X2 U2 ( .A(i5[1]), .B(n86), .C(i6[1]), .Y(n31) );
  INVX2 U3 ( .A(i5[0]), .Y(n62) );
  NOR3X4 U4 ( .A(n31), .B(n74), .C(n71), .Y(r1[1]) );
  NAND3X2TH U5 ( .A(n95), .B(n94), .C(n92), .Y(n25) );
  NOR2X4TH U6 ( .A(n53), .B(n65), .Y(r5[1]) );
  OR2XLTH U8 ( .A(n69), .B(n72), .Y(n50) );
  INVX2 U9 ( .A(i3[0]), .Y(n68) );
  OR2X2 U10 ( .A(n78), .B(n74), .Y(n54) );
  NOR2X2 U11 ( .A(n50), .B(n29), .Y(r1[3]) );
  CLKINVX1TH U12 ( .A(i1[0]), .Y(n79) );
  NAND3X2 U13 ( .A(i5[0]), .B(i4[0]), .C(i6[0]), .Y(n32) );
  NOR2X2 U14 ( .A(n54), .B(n31), .Y(r3[1]) );
  NOR3X1TH U15 ( .A(n57), .B(n26), .C(n60), .Y(r4[2]) );
  NOR3X4 U16 ( .A(n32), .B(n75), .C(n68), .Y(r1[0]) );
  NOR2X4 U17 ( .A(n51), .B(n79), .Y(r2[0]) );
  CLKINVX1TH U18 ( .A(n86), .Y(n65) );
  NAND3X3TH U19 ( .A(n87), .B(n81), .C(i2[2]), .Y(n26) );
  INVXLTH U20 ( .A(i6[1]), .Y(n58) );
  NOR3X4TH U21 ( .A(n29), .B(n76), .C(n72), .Y(r3[3]) );
  INVX2TH U22 ( .A(i2[0]), .Y(n75) );
  NOR2X6TH U23 ( .A(n52), .B(n28), .Y(r6[0]) );
  OR2XLTH U24 ( .A(n32), .B(n68), .Y(n51) );
  OR2X1TH U25 ( .A(n66), .B(n62), .Y(n52) );
  OR2XLTH U26 ( .A(n27), .B(n58), .Y(n53) );
  NOR3X1TH U27 ( .A(n57), .B(n26), .C(n67), .Y(r5[2]) );
  INVX1TH U28 ( .A(i4[0]), .Y(n66) );
  NOR3X1TH U30 ( .A(n29), .B(n76), .C(n69), .Y(r2[3]) );
  INVXLTH U31 ( .A(i1[1]), .Y(n78) );
  INVXLTH U33 ( .A(i2[2]), .Y(n73) );
  CLKINVX1TH U35 ( .A(n87), .Y(n70) );
  CLKINVX1TH U36 ( .A(i3[1]), .Y(n71) );
  NOR3X4TH U37 ( .A(n59), .B(n28), .C(n62), .Y(r4[0]) );
  NOR3X4TH U38 ( .A(n31), .B(n78), .C(n71), .Y(r2[1]) );
  OR2XLTH U39 ( .A(n73), .B(n30), .Y(n55) );
  NOR2X8 U42 ( .A(n55), .B(n70), .Y(r1[2]) );
  INVXLTH U43 ( .A(n96), .Y(n56) );
  INVXLTH U44 ( .A(n94), .Y(n76) );
  NAND3X2TH U45 ( .A(n97), .B(n93), .C(n96), .Y(n29) );
  INVXLTH U46 ( .A(n92), .Y(n69) );
  INVXLTH U47 ( .A(n95), .Y(n72) );
  INVXLTH U48 ( .A(n93), .Y(n64) );
  INVXLTH U49 ( .A(n97), .Y(n63) );
  CLKINVX1TH U51 ( .A(i6[0]), .Y(n59) );
  NOR3X1TH U52 ( .A(n56), .B(n25), .C(n63), .Y(r4[3]) );
  INVXLTH U53 ( .A(i2[1]), .Y(n74) );
  NAND3X4 U54 ( .A(i2[0]), .B(i1[0]), .C(i3[0]), .Y(n28) );
  NOR3X2 U55 ( .A(n58), .B(n27), .C(n61), .Y(r4[1]) );
  NOR3X1 U56 ( .A(n30), .B(n70), .C(n77), .Y(r2[2]) );
  INVXLTH U57 ( .A(n81), .Y(n77) );
  INVXLTH U58 ( .A(n83), .Y(n57) );
  INVXLTH U59 ( .A(i5[1]), .Y(n61) );
  INVXLTH U60 ( .A(n85), .Y(n60) );
  INVXLTH U61 ( .A(n84), .Y(n67) );
  NOR3X4TH U62 ( .A(n32), .B(n79), .C(n75), .Y(r3[0]) );
  AND3X8 U7 ( .A(n85), .B(n84), .C(n83), .Y(n80) );
  CLKINVX40 U29 ( .A(n80), .Y(n30) );
  CLKBUFX40 U32 ( .A(n88), .Y(n81) );
  INVXLTH U40 ( .A(n81), .Y(n82) );
  DLY1X1TH U41 ( .A(i6[2]), .Y(n83) );
  DLY1X1TH U50 ( .A(i4[2]), .Y(n84) );
  DLY1X1TH U63 ( .A(i5[2]), .Y(n85) );
  DLY1X1TH U64 ( .A(i4[1]), .Y(n86) );
  DLY1X1TH U65 ( .A(i3[2]), .Y(n87) );
  DLY1X1TH U66 ( .A(i1[2]), .Y(n88) );
  INVXLTH U67 ( .A(i2[2]), .Y(n89) );
  INVXLTH U68 ( .A(i5[1]), .Y(n90) );
  DLY1X1TH U69 ( .A(n64), .Y(n91) );
  DLY1X1TH U70 ( .A(i3[3]), .Y(n92) );
  DLY1X1TH U71 ( .A(i4[3]), .Y(n93) );
  DLY1X1TH U72 ( .A(i1[3]), .Y(n94) );
  DLY1X1TH U73 ( .A(i2[3]), .Y(n95) );
  DLY1X1TH U74 ( .A(i6[3]), .Y(n96) );
  DLY1X1TH U75 ( .A(i5[3]), .Y(n97) );
  OR3X8 U76 ( .A(n82), .B(n30), .C(n89), .Y(n98) );
  CLKINVX40 U77 ( .A(n98), .Y(r3[2]) );
  OR3X8 U78 ( .A(n59), .B(n28), .C(n66), .Y(n99) );
  CLKINVX40 U79 ( .A(n99), .Y(r5[0]) );
  OR3X8 U80 ( .A(n90), .B(n27), .C(n65), .Y(n100) );
  CLKINVX40 U81 ( .A(n100), .Y(r6[1]) );
  NOR3BX4 U82 ( .AN(n96), .B(n25), .C(n91), .Y(r5[3]) );
  NOR3BX4 U83 ( .AN(n97), .B(n25), .C(n91), .Y(r6[3]) );
endmodule


module sign_xor_3 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n6, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26;

  XOR2X1 U1 ( .A(n25), .B(n21), .Y(out4) );
  XOR2X3 U3 ( .A(n22), .B(in2), .Y(n6) );
  INVXLTH U4 ( .A(n4), .Y(n17) );
  XOR2XLTH U5 ( .A(in2), .B(n21), .Y(out2) );
  NAND2XLTH U6 ( .A(n18), .B(n19), .Y(out1) );
  NAND2XLTH U7 ( .A(n16), .B(n4), .Y(n19) );
  NAND2XLTH U8 ( .A(n2), .B(n17), .Y(n18) );
  INVXLTH U9 ( .A(n2), .Y(n16) );
  XNOR2X4 U10 ( .A(n3), .B(n26), .Y(n4) );
  XOR2X1TH U11 ( .A(n24), .B(n21), .Y(out3) );
  XOR2X3TH U12 ( .A(in6), .B(in5), .Y(n5) );
  XOR2XLTH U13 ( .A(in5), .B(n21), .Y(out5) );
  XNOR2X4 U14 ( .A(n2), .B(n3), .Y(n1) );
  XOR2X4 U15 ( .A(n25), .B(n5), .Y(n3) );
  XNOR2X4 U16 ( .A(n26), .B(n6), .Y(n2) );
  XNOR2X1 U2 ( .A(in6), .B(n20), .Y(out6) );
  CLKINVX40 U17 ( .A(n1), .Y(n20) );
  CLKINVX40 U18 ( .A(n20), .Y(n21) );
  DLY1X1TH U19 ( .A(in3), .Y(n22) );
  INVXLTH U20 ( .A(n22), .Y(n23) );
  INVXLTH U21 ( .A(n23), .Y(n24) );
  DLY1X1TH U22 ( .A(in4), .Y(n25) );
  DLY1X1TH U23 ( .A(in1), .Y(n26) );
endmodule


module all6_3 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88;

  NOR3X1 U50 ( .A(n30), .B(n67), .C(n59), .Y(r2[2]) );
  sign_xor_3 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR2X6 U1 ( .A(n45), .B(n28), .Y(r4[0]) );
  NOR3X4 U2 ( .A(n53), .B(n28), .C(n57), .Y(r6[0]) );
  OR2XLTH U4 ( .A(n53), .B(n49), .Y(n45) );
  NAND3X2 U5 ( .A(i6[1]), .B(n79), .C(n78), .Y(n31) );
  CLKINVX1TH U6 ( .A(i6[0]), .Y(n49) );
  CLKINVX1 U7 ( .A(n85), .Y(n53) );
  NOR3X2TH U8 ( .A(n29), .B(n66), .C(n62), .Y(r3[3]) );
  NOR3X4 U9 ( .A(n31), .B(n64), .C(n60), .Y(r1[1]) );
  NOR3X4 U10 ( .A(n32), .B(n65), .C(n61), .Y(r1[0]) );
  INVX1 U11 ( .A(n87), .Y(n61) );
  INVXL U12 ( .A(n81), .Y(n69) );
  INVX2 U13 ( .A(n88), .Y(n65) );
  NOR3X4TH U14 ( .A(n47), .B(n27), .C(n55), .Y(r5[1]) );
  NOR3X4 U15 ( .A(n49), .B(n28), .C(n57), .Y(r5[0]) );
  NAND3X2 U16 ( .A(i2[1]), .B(n80), .C(n84), .Y(n27) );
  NAND3X2TH U17 ( .A(i3[2]), .B(n77), .C(n72), .Y(n26) );
  NOR3X1TH U18 ( .A(n46), .B(n26), .C(n54), .Y(r5[2]) );
  NOR3X1TH U19 ( .A(n51), .B(n26), .C(n54), .Y(r6[2]) );
  NOR3X1TH U20 ( .A(n48), .B(n25), .C(n50), .Y(r4[3]) );
  NAND3X2TH U21 ( .A(n82), .B(n76), .C(n73), .Y(n29) );
  INVXLTH U22 ( .A(i3[3]), .Y(n58) );
  INVXLTH U23 ( .A(n75), .Y(n54) );
  INVXLTH U24 ( .A(n79), .Y(n55) );
  INVXLTH U25 ( .A(n83), .Y(n51) );
  INVXLTH U26 ( .A(n82), .Y(n50) );
  NAND3X2TH U27 ( .A(i2[3]), .B(i1[3]), .C(i3[3]), .Y(n25) );
  NOR3X1TH U28 ( .A(n29), .B(n62), .C(n58), .Y(r1[3]) );
  NOR3X2TH U29 ( .A(n46), .B(n26), .C(n51), .Y(r4[2]) );
  NAND3X3TH U30 ( .A(n85), .B(n86), .C(i6[0]), .Y(n32) );
  CLKINVX1TH U31 ( .A(i6[1]), .Y(n47) );
  NOR3X4TH U32 ( .A(n31), .B(n68), .C(n60), .Y(r2[1]) );
  CLKINVX1TH U33 ( .A(n84), .Y(n60) );
  INVXLTH U34 ( .A(n78), .Y(n52) );
  NOR3X4 U35 ( .A(n47), .B(n27), .C(n52), .Y(r4[1]) );
  INVXLTH U36 ( .A(i2[3]), .Y(n62) );
  INVXLTH U37 ( .A(n73), .Y(n48) );
  NOR3X1TH U38 ( .A(n48), .B(n25), .C(n56), .Y(r5[3]) );
  INVXLTH U39 ( .A(i1[3]), .Y(n66) );
  NOR3X1TH U40 ( .A(n50), .B(n25), .C(n56), .Y(r6[3]) );
  INVXLTH U41 ( .A(n76), .Y(n56) );
  INVXLTH U42 ( .A(n74), .Y(n46) );
  NOR3X1TH U43 ( .A(n29), .B(n66), .C(n58), .Y(r2[3]) );
  CLKINVX1TH U45 ( .A(n86), .Y(n57) );
  NOR3X2 U46 ( .A(n31), .B(n68), .C(n64), .Y(r3[1]) );
  INVXLTH U47 ( .A(n77), .Y(n67) );
  INVXLTH U48 ( .A(i3[2]), .Y(n59) );
  NOR3X2 U49 ( .A(n52), .B(n27), .C(n55), .Y(r6[1]) );
  NOR3X4TH U51 ( .A(n32), .B(n69), .C(n61), .Y(r2[0]) );
  NOR3XLTH U52 ( .A(n30), .B(n67), .C(n63), .Y(r3[2]) );
  NOR3XLTH U53 ( .A(n30), .B(n63), .C(n59), .Y(r1[2]) );
  INVXLTH U54 ( .A(n80), .Y(n68) );
  INVXLTH U55 ( .A(i2[1]), .Y(n64) );
  INVXLTH U56 ( .A(n72), .Y(n63) );
  NOR3XLTH U57 ( .A(n32), .B(n69), .C(n65), .Y(r3[0]) );
  AND3X8 U3 ( .A(n88), .B(n81), .C(n87), .Y(n70) );
  CLKINVX40 U44 ( .A(n70), .Y(n28) );
  AND3X8 U58 ( .A(n83), .B(n75), .C(n74), .Y(n71) );
  CLKINVX40 U59 ( .A(n71), .Y(n30) );
  DLY1X1TH U60 ( .A(i2[2]), .Y(n72) );
  DLY1X1TH U61 ( .A(i6[3]), .Y(n73) );
  DLY1X1TH U62 ( .A(i6[2]), .Y(n74) );
  DLY1X1TH U63 ( .A(i4[2]), .Y(n75) );
  DLY1X1TH U64 ( .A(i4[3]), .Y(n76) );
  DLY1X1TH U65 ( .A(i1[2]), .Y(n77) );
  DLY1X1TH U66 ( .A(i5[1]), .Y(n78) );
  DLY1X1TH U67 ( .A(i4[1]), .Y(n79) );
  DLY1X1TH U68 ( .A(i1[1]), .Y(n80) );
  DLY1X1TH U69 ( .A(i1[0]), .Y(n81) );
  DLY1X1TH U70 ( .A(i5[3]), .Y(n82) );
  DLY1X1TH U71 ( .A(i5[2]), .Y(n83) );
  DLY1X1TH U72 ( .A(i3[1]), .Y(n84) );
  DLY1X1TH U73 ( .A(i5[0]), .Y(n85) );
  DLY1X1TH U74 ( .A(i4[0]), .Y(n86) );
  DLY1X1TH U75 ( .A(i3[0]), .Y(n87) );
  DLY1X1TH U76 ( .A(i2[0]), .Y(n88) );
endmodule


module sign_xor_2 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n4, n5, n25, n26, n27, n28, n29, n30;

  XOR2X1 U1 ( .A(in2), .B(n1), .Y(out2) );
  XOR2XL U2 ( .A(n30), .B(n1), .Y(out1) );
  XOR2XL U3 ( .A(in4), .B(n1), .Y(out4) );
  CLKXOR2X8 U4 ( .A(n2), .B(n25), .Y(n1) );
  XOR2X3 U5 ( .A(n26), .B(in2), .Y(n5) );
  XNOR2X4TH U6 ( .A(in1), .B(n5), .Y(n2) );
  XOR2X2TH U7 ( .A(in6), .B(in5), .Y(n4) );
  XOR2XLTH U8 ( .A(n28), .B(n1), .Y(out3) );
  XOR2X1TH U9 ( .A(in6), .B(n1), .Y(out6) );
  XOR2X1TH U10 ( .A(in5), .B(n1), .Y(out5) );
  XNOR2X4 U11 ( .A(in4), .B(n4), .Y(n25) );
  DLY1X1TH U12 ( .A(in3), .Y(n26) );
  INVXLTH U13 ( .A(n26), .Y(n27) );
  INVXLTH U14 ( .A(n27), .Y(n28) );
  INVXLTH U15 ( .A(in1), .Y(n29) );
  INVXLTH U16 ( .A(n29), .Y(n30) );
endmodule


module all6_2 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87;

  NAND3X2 U5 ( .A(n83), .B(n81), .C(n79), .Y(n29) );
  sign_xor_2 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X1 U1 ( .A(n49), .B(n45), .C(n53), .Y(r4[0]) );
  NOR2X4 U2 ( .A(n44), .B(n69), .Y(r3[0]) );
  NAND3X4 U3 ( .A(n76), .B(i4[1]), .C(i5[1]), .Y(n31) );
  INVX1 U4 ( .A(n77), .Y(n63) );
  BUFX3TH U7 ( .A(n28), .Y(n45) );
  NAND3X2 U8 ( .A(n86), .B(n75), .C(n71), .Y(n32) );
  NAND3X2 U9 ( .A(n85), .B(n82), .C(n80), .Y(n25) );
  NOR3X1 U10 ( .A(n48), .B(n26), .C(n51), .Y(r4[2]) );
  OR2X2TH U11 ( .A(n32), .B(n64), .Y(n44) );
  NAND3X2 U12 ( .A(i5[2]), .B(i4[2]), .C(i6[2]), .Y(n30) );
  INVX2 U13 ( .A(n86), .Y(n53) );
  INVX1 U14 ( .A(i1[0]), .Y(n69) );
  INVX1 U15 ( .A(n84), .Y(n64) );
  NOR3X1TH U16 ( .A(n30), .B(n67), .C(n62), .Y(r3[2]) );
  NOR3X4TH U17 ( .A(n31), .B(n63), .C(n59), .Y(r1[1]) );
  INVXLTH U18 ( .A(i5[2]), .Y(n51) );
  INVXLTH U19 ( .A(n72), .Y(n61) );
  INVXLTH U20 ( .A(n74), .Y(n60) );
  NOR3X2 U21 ( .A(n32), .B(n64), .C(n60), .Y(r1[0]) );
  INVX2TH U22 ( .A(n85), .Y(n65) );
  INVXLTH U23 ( .A(n82), .Y(n66) );
  NOR3X1TH U24 ( .A(n47), .B(n25), .C(n50), .Y(r4[3]) );
  INVXLTH U25 ( .A(n73), .Y(n62) );
  NOR3X1TH U26 ( .A(n30), .B(n62), .C(n61), .Y(r1[2]) );
  NOR3X1TH U27 ( .A(n47), .B(n25), .C(n54), .Y(r5[3]) );
  INVXLTH U28 ( .A(n80), .Y(n58) );
  NAND3X4TH U29 ( .A(n77), .B(i1[1]), .C(i3[1]), .Y(n27) );
  NOR3X1TH U30 ( .A(n29), .B(n66), .C(n58), .Y(r2[3]) );
  INVXLTH U31 ( .A(i1[2]), .Y(n67) );
  INVXLTH U32 ( .A(i1[1]), .Y(n68) );
  CLKINVX1TH U33 ( .A(i3[1]), .Y(n59) );
  NOR3X4TH U34 ( .A(n51), .B(n26), .C(n56), .Y(r6[2]) );
  NOR3X1TH U35 ( .A(n50), .B(n25), .C(n54), .Y(r6[3]) );
  NOR3X4TH U36 ( .A(n46), .B(n27), .C(n55), .Y(r5[1]) );
  NOR3XLTH U37 ( .A(n48), .B(n26), .C(n56), .Y(r5[2]) );
  NAND3X2TH U38 ( .A(i1[0]), .B(n84), .C(n74), .Y(n28) );
  NOR3X4TH U39 ( .A(n31), .B(n68), .C(n59), .Y(r2[1]) );
  NOR3X4TH U40 ( .A(n32), .B(n69), .C(n60), .Y(r2[0]) );
  NOR3X2 U41 ( .A(n46), .B(n27), .C(n52), .Y(r4[1]) );
  NOR3X2 U42 ( .A(n52), .B(n27), .C(n55), .Y(r6[1]) );
  NOR3X2 U43 ( .A(n31), .B(n68), .C(n63), .Y(r3[1]) );
  INVXLTH U44 ( .A(i4[1]), .Y(n55) );
  NOR3XLTH U45 ( .A(n30), .B(n67), .C(n61), .Y(r2[2]) );
  NOR3X1TH U46 ( .A(n29), .B(n65), .C(n58), .Y(r1[3]) );
  NOR3X1TH U47 ( .A(n29), .B(n66), .C(n65), .Y(r3[3]) );
  INVXLTH U48 ( .A(n71), .Y(n49) );
  INVXLTH U49 ( .A(n76), .Y(n46) );
  INVXLTH U50 ( .A(i6[2]), .Y(n48) );
  INVXLTH U51 ( .A(n79), .Y(n47) );
  INVXLTH U52 ( .A(i5[1]), .Y(n52) );
  INVXLTH U53 ( .A(n83), .Y(n50) );
  INVXLTH U54 ( .A(i4[2]), .Y(n56) );
  INVXLTH U55 ( .A(n81), .Y(n54) );
  CLKINVX1TH U56 ( .A(n75), .Y(n57) );
  NOR3X4 U57 ( .A(n53), .B(n45), .C(n57), .Y(r6[0]) );
  AND3X8 U6 ( .A(i1[2]), .B(n73), .C(n72), .Y(n70) );
  CLKINVX40 U58 ( .A(n70), .Y(n26) );
  DLY1X1TH U59 ( .A(i6[0]), .Y(n71) );
  DLY1X1TH U60 ( .A(i3[2]), .Y(n72) );
  DLY1X1TH U61 ( .A(i2[2]), .Y(n73) );
  DLY1X1TH U62 ( .A(i3[0]), .Y(n74) );
  DLY1X1TH U63 ( .A(i4[0]), .Y(n75) );
  DLY1X1TH U64 ( .A(i6[1]), .Y(n76) );
  DLY1X1TH U65 ( .A(i2[1]), .Y(n77) );
  DLY1X1TH U66 ( .A(n49), .Y(n78) );
  DLY1X1TH U67 ( .A(i6[3]), .Y(n79) );
  DLY1X1TH U68 ( .A(i3[3]), .Y(n80) );
  DLY1X1TH U69 ( .A(i4[3]), .Y(n81) );
  DLY1X1TH U70 ( .A(i1[3]), .Y(n82) );
  DLY1X1TH U71 ( .A(i5[3]), .Y(n83) );
  DLY1X1TH U72 ( .A(i2[0]), .Y(n84) );
  DLY1X1TH U73 ( .A(i2[3]), .Y(n85) );
  DLY1X1TH U74 ( .A(i5[0]), .Y(n86) );
  OR3X8 U75 ( .A(n78), .B(n45), .C(n57), .Y(n87) );
  CLKINVX40 U76 ( .A(n87), .Y(r5[0]) );
endmodule


module sign_xor_1 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n2, n3, n4, n5, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33;

  CLKNAND2X2 U1 ( .A(in1), .B(n21), .Y(n22) );
  NAND2XLTH U2 ( .A(n20), .B(n1), .Y(n23) );
  NAND2X2 U3 ( .A(n22), .B(n23), .Y(out1) );
  INVXLTH U4 ( .A(in1), .Y(n20) );
  CLKINVX3 U5 ( .A(n1), .Y(n21) );
  BUFX6 U7 ( .A(in6), .Y(n24) );
  XOR2X4 U8 ( .A(n24), .B(in5), .Y(n4) );
  XOR2X1TH U9 ( .A(in5), .B(n1), .Y(out5) );
  NAND2X1 U10 ( .A(n2), .B(n3), .Y(n27) );
  INVX10 U11 ( .A(n2), .Y(n25) );
  XNOR2X4 U12 ( .A(in1), .B(n5), .Y(n2) );
  CLKNAND2X8 U13 ( .A(n27), .B(n28), .Y(n1) );
  XOR2X1 U14 ( .A(in3), .B(in2), .Y(n5) );
  XOR2X4 U15 ( .A(n31), .B(n4), .Y(n3) );
  XOR2XL U16 ( .A(n24), .B(n1), .Y(out6) );
  XOR2X1 U18 ( .A(n33), .B(n1), .Y(out4) );
  CLKNAND2X4 U19 ( .A(n25), .B(n26), .Y(n28) );
  INVX1TH U20 ( .A(n3), .Y(n26) );
  XNOR2X1 U6 ( .A(n29), .B(n1), .Y(out2) );
  CLKINVX40 U17 ( .A(in2), .Y(n29) );
  XNOR2X1 U21 ( .A(n30), .B(n1), .Y(out3) );
  CLKINVX40 U22 ( .A(in3), .Y(n30) );
  DLY1X1TH U23 ( .A(in4), .Y(n31) );
  INVXLTH U24 ( .A(n31), .Y(n32) );
  INVXLTH U25 ( .A(n32), .Y(n33) );
endmodule


module all6_1 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93;

  NOR3X1 U41 ( .A(n51), .B(n25), .C(n55), .Y(r4[3]) );
  sign_xor_1 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X4 U1 ( .A(n57), .B(n27), .C(n62), .Y(r6[1]) );
  NOR3X4 U2 ( .A(n32), .B(n74), .C(n66), .Y(r2[0]) );
  NOR3XL U3 ( .A(n32), .B(n69), .C(n66), .Y(r1[0]) );
  NAND3X2 U4 ( .A(n86), .B(n88), .C(n82), .Y(n31) );
  NOR3X4 U5 ( .A(n54), .B(n28), .C(n56), .Y(r4[0]) );
  AND2XLTH U6 ( .A(n77), .B(n78), .Y(n47) );
  NOR2X4 U7 ( .A(n64), .B(n68), .Y(n48) );
  NOR2X2 U8 ( .A(n49), .B(n31), .Y(r1[1]) );
  INVX2 U9 ( .A(n48), .Y(n49) );
  NAND2X4 U10 ( .A(i1[0]), .B(n47), .Y(n28) );
  NOR3X4 U13 ( .A(n53), .B(n27), .C(n62), .Y(r5[1]) );
  NAND3X2 U14 ( .A(i2[1]), .B(i1[1]), .C(i3[1]), .Y(n27) );
  NOR3X4TH U15 ( .A(n32), .B(n74), .C(n69), .Y(r3[0]) );
  NAND3X2 U16 ( .A(n87), .B(n84), .C(n83), .Y(n30) );
  NOR3X2 U17 ( .A(n31), .B(n73), .C(n64), .Y(r2[1]) );
  INVX2TH U18 ( .A(i4[0]), .Y(n60) );
  INVXLTH U19 ( .A(i1[1]), .Y(n73) );
  CLKINVX1TH U20 ( .A(n77), .Y(n66) );
  NOR3X4TH U21 ( .A(n29), .B(n70), .C(n65), .Y(r1[3]) );
  NOR3X1TH U22 ( .A(n52), .B(n26), .C(n61), .Y(r5[2]) );
  INVX2TH U23 ( .A(n91), .Y(n56) );
  NOR3X1 U24 ( .A(n31), .B(n73), .C(n68), .Y(r3[1]) );
  CLKINVX1TH U25 ( .A(n88), .Y(n62) );
  INVX1TH U27 ( .A(n90), .Y(n54) );
  INVX2TH U28 ( .A(n89), .Y(n63) );
  NOR3X4TH U29 ( .A(n52), .B(n26), .C(n58), .Y(r4[2]) );
  OR2XLTH U30 ( .A(n30), .B(n63), .Y(n50) );
  CLKINVX1TH U31 ( .A(n78), .Y(n69) );
  NOR3XLTH U33 ( .A(n30), .B(n72), .C(n67), .Y(r3[2]) );
  NOR3X1TH U34 ( .A(n30), .B(n72), .C(n63), .Y(r2[2]) );
  NOR3X1TH U35 ( .A(n58), .B(n26), .C(n61), .Y(r6[2]) );
  NOR3X1TH U36 ( .A(n51), .B(n25), .C(n59), .Y(r5[3]) );
  NOR3X1TH U37 ( .A(n29), .B(n71), .C(n70), .Y(r3[3]) );
  NOR3X1TH U38 ( .A(n29), .B(n71), .C(n65), .Y(r2[3]) );
  INVXLTH U39 ( .A(n80), .Y(n59) );
  NAND3X2TH U40 ( .A(i2[3]), .B(i1[3]), .C(i3[3]), .Y(n25) );
  INVXLTH U42 ( .A(n85), .Y(n55) );
  INVXLTH U43 ( .A(n79), .Y(n51) );
  INVXLTH U44 ( .A(i1[3]), .Y(n71) );
  INVXLTH U45 ( .A(i2[3]), .Y(n70) );
  NAND3X2TH U46 ( .A(n85), .B(n80), .C(n79), .Y(n29) );
  INVXLTH U47 ( .A(i3[3]), .Y(n65) );
  NOR3X1TH U48 ( .A(n55), .B(n25), .C(n59), .Y(r6[3]) );
  INVXLTH U49 ( .A(n82), .Y(n53) );
  INVXLTH U50 ( .A(n81), .Y(n72) );
  INVXLTH U51 ( .A(i2[1]), .Y(n68) );
  INVXLTH U52 ( .A(n86), .Y(n57) );
  INVXLTH U53 ( .A(n83), .Y(n52) );
  INVXLTH U54 ( .A(n84), .Y(n61) );
  INVXLTH U55 ( .A(i2[2]), .Y(n67) );
  INVX2 U56 ( .A(i1[0]), .Y(n74) );
  NOR3X2 U57 ( .A(n53), .B(n27), .C(n57), .Y(r4[1]) );
  NAND3X4 U58 ( .A(n91), .B(i4[0]), .C(n90), .Y(n32) );
  INVXLTH U59 ( .A(n87), .Y(n58) );
  INVXLTH U60 ( .A(i3[1]), .Y(n64) );
  OR3X8 U11 ( .A(n56), .B(n28), .C(n60), .Y(n75) );
  CLKINVX40 U12 ( .A(n75), .Y(r6[0]) );
  AND3X8 U26 ( .A(i2[2]), .B(n81), .C(n89), .Y(n76) );
  CLKINVX40 U32 ( .A(n76), .Y(n26) );
  DLY1X1TH U61 ( .A(i3[0]), .Y(n77) );
  DLY1X1TH U62 ( .A(i2[0]), .Y(n78) );
  DLY1X1TH U63 ( .A(i6[3]), .Y(n79) );
  DLY1X1TH U64 ( .A(i4[3]), .Y(n80) );
  DLY1X1TH U65 ( .A(i1[2]), .Y(n81) );
  DLY1X1TH U66 ( .A(i6[1]), .Y(n82) );
  DLY1X1TH U67 ( .A(i6[2]), .Y(n83) );
  DLY1X1TH U68 ( .A(i4[2]), .Y(n84) );
  DLY1X1TH U69 ( .A(i5[3]), .Y(n85) );
  DLY1X1TH U70 ( .A(i5[1]), .Y(n86) );
  DLY1X1TH U71 ( .A(i5[2]), .Y(n87) );
  DLY1X1TH U72 ( .A(i4[1]), .Y(n88) );
  DLY1X1TH U73 ( .A(i3[2]), .Y(n89) );
  DLY1X1TH U74 ( .A(i6[0]), .Y(n90) );
  DLY1X1TH U75 ( .A(i5[0]), .Y(n91) );
  OR2X8 U76 ( .A(n50), .B(n67), .Y(n92) );
  CLKINVX40 U77 ( .A(n92), .Y(r1[2]) );
  OR3X8 U78 ( .A(n54), .B(n28), .C(n60), .Y(n93) );
  CLKINVX40 U79 ( .A(n93), .Y(r5[0]) );
endmodule


module sign_xor_0 ( out1, out2, out3, out4, out5, out6, in1, in2, in3, in4, 
        in5, in6 );
  input in1, in2, in3, in4, in5, in6;
  output out1, out2, out3, out4, out5, out6;
  wire   n1, n3, n4, n5, n20, n21, n22, n23, n24, n25;

  XOR2X1 U1 ( .A(in1), .B(n1), .Y(out1) );
  XOR2X1 U2 ( .A(in2), .B(n1), .Y(out2) );
  XOR2X1 U3 ( .A(in4), .B(n1), .Y(out4) );
  NAND2X2 U4 ( .A(in3), .B(n21), .Y(n22) );
  NAND2XL U5 ( .A(n20), .B(n1), .Y(n23) );
  NAND2X2 U6 ( .A(n22), .B(n23), .Y(out3) );
  INVXLTH U7 ( .A(in3), .Y(n20) );
  INVXL U8 ( .A(n1), .Y(n21) );
  CLKXOR2X12 U9 ( .A(n24), .B(n3), .Y(n1) );
  XOR2X1 U10 ( .A(in6), .B(in5), .Y(n4) );
  XOR2XL U12 ( .A(in6), .B(n1), .Y(out6) );
  XOR2X2TH U13 ( .A(in4), .B(n4), .Y(n3) );
  XOR2X3TH U14 ( .A(in3), .B(in2), .Y(n5) );
  XOR2X4 U15 ( .A(in1), .B(n5), .Y(n24) );
  XNOR2X1 U11 ( .A(n25), .B(n1), .Y(out5) );
  CLKINVX40 U16 ( .A(in5), .Y(n25) );
endmodule


module all6_0 ( r1, r2, r3, r4, r5, r6, i1, i2, i3, i4, i5, i6 );
  output [4:0] r1;
  output [4:0] r2;
  output [4:0] r3;
  output [4:0] r4;
  output [4:0] r5;
  output [4:0] r6;
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n44, n45, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88;

  sign_xor_0 sign_xor_1 ( .out1(r1[4]), .out2(r2[4]), .out3(r3[4]), .out4(
        r4[4]), .out5(r5[4]), .out6(r6[4]), .in1(i1[4]), .in2(i2[4]), .in3(
        i3[4]), .in4(i4[4]), .in5(i5[4]), .in6(i6[4]) );
  NOR3X1 U1 ( .A(n30), .B(n67), .C(n60), .Y(r2[2]) );
  INVX2 U4 ( .A(i2[2]), .Y(n64) );
  NOR3X1 U6 ( .A(n49), .B(n28), .C(n57), .Y(r5[0]) );
  NOR3X4 U7 ( .A(n50), .B(n27), .C(n54), .Y(r4[1]) );
  NAND3X2 U8 ( .A(i5[1]), .B(i4[1]), .C(n76), .Y(n31) );
  NAND3X2 U9 ( .A(n79), .B(n78), .C(n77), .Y(n32) );
  INVXL U10 ( .A(n74), .Y(n62) );
  OR2XLTH U11 ( .A(n57), .B(n53), .Y(n45) );
  NOR3X1TH U12 ( .A(n30), .B(n64), .C(n60), .Y(r1[2]) );
  NOR3X2TH U13 ( .A(n32), .B(n65), .C(n61), .Y(r1[0]) );
  NOR3X1TH U14 ( .A(n47), .B(n26), .C(n52), .Y(r4[2]) );
  NOR3X4 U16 ( .A(n30), .B(n67), .C(n64), .Y(r3[2]) );
  NAND3X2TH U17 ( .A(i5[2]), .B(i4[2]), .C(i6[2]), .Y(n30) );
  INVXLTH U18 ( .A(i1[2]), .Y(n67) );
  NOR3X4 U19 ( .A(n49), .B(n28), .C(n53), .Y(r4[0]) );
  NOR3X1TH U20 ( .A(n29), .B(n69), .C(n63), .Y(r3[3]) );
  INVXLTH U21 ( .A(i4[2]), .Y(n56) );
  INVX1TH U22 ( .A(n79), .Y(n53) );
  NOR3XLTH U23 ( .A(n52), .B(n26), .C(n56), .Y(r6[2]) );
  NOR3X4TH U24 ( .A(n31), .B(n66), .C(n62), .Y(r1[1]) );
  OR2XLTH U25 ( .A(n70), .B(n65), .Y(n44) );
  NAND3X4 U26 ( .A(n80), .B(i1[2]), .C(i2[2]), .Y(n26) );
  NOR3X2TH U27 ( .A(n29), .B(n69), .C(n59), .Y(r2[3]) );
  NOR3X1TH U28 ( .A(n48), .B(n25), .C(n51), .Y(r4[3]) );
  INVXLTH U29 ( .A(i4[3]), .Y(n55) );
  NAND3X2TH U30 ( .A(n85), .B(n84), .C(n83), .Y(n25) );
  INVXLTH U31 ( .A(i5[3]), .Y(n51) );
  INVXLTH U32 ( .A(i6[3]), .Y(n48) );
  INVXLTH U33 ( .A(n84), .Y(n69) );
  NAND3X2TH U34 ( .A(i5[3]), .B(i4[3]), .C(i6[3]), .Y(n29) );
  INVXLTH U35 ( .A(n83), .Y(n59) );
  INVXLTH U36 ( .A(n85), .Y(n63) );
  NOR3X1TH U37 ( .A(n51), .B(n25), .C(n55), .Y(r6[3]) );
  NOR3X1TH U38 ( .A(n48), .B(n25), .C(n55), .Y(r5[3]) );
  NAND3X2TH U39 ( .A(i1[1]), .B(n75), .C(n74), .Y(n27) );
  NOR3X1TH U40 ( .A(n29), .B(n63), .C(n59), .Y(r1[3]) );
  INVXLTH U41 ( .A(n75), .Y(n66) );
  INVXLTH U43 ( .A(i2[0]), .Y(n65) );
  INVXLTH U44 ( .A(i3[0]), .Y(n61) );
  NOR3X2 U46 ( .A(n54), .B(n27), .C(n58), .Y(r6[1]) );
  INVXL U48 ( .A(n78), .Y(n57) );
  INVXLTH U49 ( .A(n73), .Y(n70) );
  NOR3X2 U50 ( .A(n31), .B(n81), .C(n66), .Y(r3[1]) );
  INVXLTH U51 ( .A(n76), .Y(n50) );
  INVXLTH U52 ( .A(i6[2]), .Y(n47) );
  INVXLTH U53 ( .A(i5[2]), .Y(n52) );
  INVXLTH U54 ( .A(n77), .Y(n49) );
  INVXLTH U55 ( .A(i5[1]), .Y(n54) );
  NOR3X2 U56 ( .A(n50), .B(n27), .C(n58), .Y(r5[1]) );
  INVXLTH U57 ( .A(i1[1]), .Y(n68) );
  INVXLTH U58 ( .A(i4[1]), .Y(n58) );
  INVXLTH U59 ( .A(n80), .Y(n60) );
  NAND3BX4 U2 ( .AN(n32), .B(n73), .C(i3[0]), .Y(n71) );
  CLKINVX40 U3 ( .A(n71), .Y(r2[0]) );
  AND3X8 U5 ( .A(i2[0]), .B(i3[0]), .C(n73), .Y(n72) );
  CLKINVX40 U15 ( .A(n72), .Y(n28) );
  DLY1X1TH U42 ( .A(i1[0]), .Y(n73) );
  DLY1X1TH U45 ( .A(i3[1]), .Y(n74) );
  DLY1X1TH U47 ( .A(i2[1]), .Y(n75) );
  DLY1X1TH U60 ( .A(i6[1]), .Y(n76) );
  DLY1X1TH U61 ( .A(i6[0]), .Y(n77) );
  DLY1X1TH U62 ( .A(i4[0]), .Y(n78) );
  DLY1X1TH U63 ( .A(i5[0]), .Y(n79) );
  DLY1X1TH U64 ( .A(i3[2]), .Y(n80) );
  INVXLTH U65 ( .A(i1[1]), .Y(n81) );
  DLY1X1TH U66 ( .A(n62), .Y(n82) );
  DLY1X1TH U67 ( .A(i3[3]), .Y(n83) );
  DLY1X1TH U68 ( .A(i1[3]), .Y(n84) );
  DLY1X1TH U69 ( .A(i2[3]), .Y(n85) );
  OR3X8 U70 ( .A(n82), .B(n68), .C(n31), .Y(n86) );
  CLKINVX40 U71 ( .A(n86), .Y(r2[1]) );
  NOR3BX4 U72 ( .AN(i6[2]), .B(n26), .C(n56), .Y(r5[2]) );
  OR2X8 U73 ( .A(n45), .B(n28), .Y(n87) );
  CLKINVX40 U74 ( .A(n87), .Y(r6[0]) );
  OR2X8 U75 ( .A(n44), .B(n32), .Y(n88) );
  CLKINVX40 U76 ( .A(n88), .Y(r3[0]) );
endmodule


module sm_tc_191 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n19, n20, n23;

  XNOR2X1 U2 ( .A(n20), .B(n8), .Y(n5) );
  INVX12 U3 ( .A(in[4]), .Y(n19) );
  AOI31X1 U4 ( .A0(n3), .A1(n4), .A2(n5), .B0(n19), .Y(out[4]) );
  INVX2 U5 ( .A(in[2]), .Y(n20) );
  NOR2X6 U7 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI2BB2X2 U8 ( .B0(n19), .B1(n4), .A0N(n23), .A1N(n19), .Y(out[3]) );
  AO21XL U9 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  XNOR2X2TH U10 ( .A(n7), .B(n23), .Y(n4) );
  NAND2XLTH U11 ( .A(n8), .B(n20), .Y(n7) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX1TH U14 ( .A(in[0]), .Y(out[0]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX40 U6 ( .A(in[3]), .Y(n23) );
  AO2B2X4 U12 ( .B0(in[1]), .B1(n19), .A0(in[4]), .A1N(n6), .Y(out[1]) );
  OAI2B2X2 U17 ( .A1N(in[4]), .A0(n5), .B0(in[4]), .B1(n20), .Y(out[2]) );
endmodule


module sm_tc_190 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n19, n20, n21, n22, n26, n27;

  NOR2X4 U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U3 ( .A(in[2]), .Y(n27) );
  XNOR2X2 U4 ( .A(n27), .B(n8), .Y(n5) );
  AO21XLTH U5 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2X2 U6 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n26), .Y(out[1]) );
  BUFX2TH U7 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X1TH U8 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  NAND2X1TH U9 ( .A(n8), .B(n27), .Y(n7) );
  OAI22XL U10 ( .A0(in[4]), .A1(n27), .B0(n26), .B1(n5), .Y(out[2]) );
  INVX2TH U11 ( .A(n7), .Y(n19) );
  CLKNAND2X2TH U12 ( .A(n7), .B(in[3]), .Y(n21) );
  CLKNAND2X4 U13 ( .A(n19), .B(n20), .Y(n22) );
  CLKNAND2X8 U14 ( .A(n21), .B(n22), .Y(n4) );
  INVX1 U15 ( .A(in[3]), .Y(n20) );
  AOI31X4 U16 ( .A0(n3), .A1(n4), .A2(n5), .B0(n26), .Y(out[5]) );
  INVX3TH U17 ( .A(in[4]), .Y(n26) );
  CLKBUFX1TH U18 ( .A(out[5]), .Y(out[6]) );
  CLKBUFX1TH U19 ( .A(out[5]), .Y(out[4]) );
  NOR2BXLTH U20 ( .AN(n6), .B(in[0]), .Y(n3) );
endmodule


module sm_tc_189 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n21, n25, n26;

  NOR2X2TH U2 ( .A(in[1]), .B(out[0]), .Y(n8) );
  INVX2TH U3 ( .A(in[2]), .Y(n25) );
  OAI22XLTH U4 ( .A0(in[4]), .A1(n25), .B0(n26), .B1(n21), .Y(out[2]) );
  AO21X4 U5 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NAND2XLTH U6 ( .A(n8), .B(n25), .Y(n7) );
  XNOR2X4 U7 ( .A(n25), .B(n8), .Y(n5) );
  BUFX6 U8 ( .A(n5), .Y(n21) );
  BUFX12 U9 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X1TH U10 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n26), .Y(out[1]) );
  AOI31X4TH U11 ( .A0(n3), .A1(n4), .A2(n21), .B0(n26), .Y(out[4]) );
  NOR2BXLTH U12 ( .AN(n6), .B(out[0]), .Y(n3) );
  INVX3TH U13 ( .A(in[4]), .Y(n26) );
  XNOR2X4 U14 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X1TH U17 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
endmodule


module sm_tc_188 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  OAI2BB2X1TH U2 ( .B0(n21), .B1(n6), .A0N(in[1]), .A1N(n21), .Y(out[1]) );
  CLKBUFX1TH U3 ( .A(in[0]), .Y(out[0]) );
  OAI22X1TH U4 ( .A0(in[4]), .A1(n22), .B0(n21), .B1(n5), .Y(out[2]) );
  NOR2X3TH U5 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X1TH U6 ( .A(n7), .B(in[3]), .Y(n4) );
  INVXLTH U7 ( .A(out[4]), .Y(n18) );
  CLKINVX2TH U8 ( .A(in[4]), .Y(n21) );
  CLKINVX1TH U9 ( .A(in[2]), .Y(n22) );
  AOI31X2TH U10 ( .A0(n3), .A1(n4), .A2(n5), .B0(n21), .Y(out[4]) );
  NOR2BXLTH U11 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U12 ( .A(n18), .Y(out[5]) );
  OAI2BB2X2TH U13 ( .B0(n21), .B1(n4), .A0N(in[3]), .A1N(n21), .Y(out[3]) );
  INVXLTH U14 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U15 ( .A(n22), .B(n8), .Y(n5) );
  NAND2XLTH U16 ( .A(n8), .B(n22), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_47_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_47_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR2X4 U1 ( .A(n6), .B(A[6]), .Y(SUM[6]) );
  NAND3X4 U3 ( .A(n3), .B(n4), .C(n5), .Y(carry[4]) );
  XOR2X3 U4 ( .A(B[6]), .B(carry[6]), .Y(n6) );
  XOR2XLTH U5 ( .A(B[3]), .B(A[3]), .Y(n2) );
  CLKXOR2X1TH U6 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2XLTH U7 ( .A(A[3]), .B(B[3]), .Y(n5) );
  XOR2X1TH U9 ( .A(n2), .B(carry[3]), .Y(SUM[3]) );
  AND2XLTH U10 ( .A(B[0]), .B(A[0]), .Y(n1) );
  AND2X8 U2 ( .A(carry[3]), .B(B[3]), .Y(n7) );
  CLKINVX40 U8 ( .A(n7), .Y(n4) );
  AND2X8 U11 ( .A(carry[3]), .B(A[3]), .Y(n8) );
  CLKINVX40 U12 ( .A(n8), .Y(n3) );
endmodule


module add_47_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_47_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX4TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR2X1 U1 ( .A(A[6]), .B(B[6]), .Y(n2) );
  CLKXOR2X8 U2 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_47_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR2X1 U1 ( .A(n2), .B(A[0]), .Y(SUM[0]) );
  CLKINVX40 U3 ( .A(B[0]), .Y(n2) );
endmodule


module add_47_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_47 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n13, n14, n15, n16, n17, n18, n19, n20, n21;

  add_47_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, n21}), .B({in2[6:3], n18, n14, n13}), .SUM(out3)
         );
  add_47_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, n20, temp2_3_, temp2_2_, 
        temp2_1_, n15}), .B(in), .SUM(out1) );
  add_47_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, n21}), .B({in3[6:3], n19, in3[1:0]}), .SUM(out2)
         );
  add_47_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, n17}), .B({temp2_6_, temp2_5_, n20, temp2_3_, 
        temp2_2_, temp2_1_, n15}), .SUM(out) );
  add_47_DW01_add_4 add_30 ( .A({in2[6:3], n18, n14, n13}), .B({in3[6:3], n19, 
        in3[1:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_47_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX2TH U1 ( .A(in2[1]), .Y(n14) );
  CLKBUFX1TH U2 ( .A(temp2_0_), .Y(n15) );
  BUFX10 U3 ( .A(in2[0]), .Y(n13) );
  CLKBUFX1TH U4 ( .A(in2[2]), .Y(n18) );
  INVXLTH U5 ( .A(n21), .Y(n16) );
  INVXLTH U6 ( .A(n16), .Y(n17) );
  BUFX2TH U13 ( .A(in3[2]), .Y(n19) );
  CLKBUFX40 U14 ( .A(temp2_4_), .Y(n20) );
  CLKBUFX40 U15 ( .A(temp1_0_), .Y(n21) );
endmodule


module tc_sm_191 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n17, n18, n19, n20, n21, n22;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n22) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n21) );
  XNOR2XLTH U7 ( .A(n21), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(in[6]), .Y(n17) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n18), .B2(
        n19), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n19) );
  INVXLTH U12 ( .A(in[5]), .Y(n18) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n20) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U16 ( .A0(n17), .A1(n12), .B0(in[6]), .B1(n22), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n17), .A1(n10), .B0(in[6]), .B1(n21), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n20), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n20), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n20), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_190 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n18, n19, n20, n21, n22, n23, n25,
         n26, n27, n28, n30;

  NAND3X2 U3 ( .A(n21), .B(n22), .C(n6), .Y(out[2]) );
  INVX2 U4 ( .A(in[6]), .Y(n23) );
  CLKINVX4 U5 ( .A(out[4]), .Y(n25) );
  OAI211XL U6 ( .A0(out[4]), .A1(n26), .B0(n5), .C0(n6), .Y(out[3]) );
  CLKINVX12 U8 ( .A(n23), .Y(out[4]) );
  NOR2XL U9 ( .A(n25), .B(n10), .Y(n18) );
  NOR2XLTH U10 ( .A(out[4]), .B(n28), .Y(n19) );
  INVXLTH U11 ( .A(n6), .Y(n20) );
  OR3X2TH U12 ( .A(n18), .B(n19), .C(n20), .Y(out[1]) );
  AOI21X8 U13 ( .A0(out[4]), .A1(n11), .B0(n12), .Y(n6) );
  OAI2B11X2TH U14 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  AOI2BB1X1TH U15 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  NOR3X1TH U16 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  XOR2XLTH U17 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n9) );
  XOR2XLTH U19 ( .A(in[0]), .B(n28), .Y(n10) );
  INVXLTH U20 ( .A(in[1]), .Y(n28) );
  INVXLTH U21 ( .A(in[3]), .Y(n26) );
  OR2XLTH U22 ( .A(out[4]), .B(n27), .Y(n22) );
  OR2XLTH U23 ( .A(n25), .B(n8), .Y(n21) );
  INVXLTH U24 ( .A(in[2]), .Y(n27) );
  NAND2BXLTH U25 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  OA21X4 U7 ( .A0(n7), .A1(n26), .B0(out[4]), .Y(n30) );
  CLKINVX40 U26 ( .A(n30), .Y(n5) );
endmodule


module tc_sm_189 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n17, n19, n20, n21, n22, n23, n24;

  BUFX6 U3 ( .A(n8), .Y(n17) );
  OAI221XL U4 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n17), .Y(out[1])
         );
  OAI221XL U5 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n17), .Y(out[2])
         );
  OAI211XL U6 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n17), .Y(out[3]) );
  CLKINVX1TH U7 ( .A(in[3]), .Y(n22) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  OAI33X4 U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n20), .B2(n21), .Y(n8) );
  OAI2BB1X4 U10 ( .A0N(n22), .A1N(n9), .B0(in[6]), .Y(n13) );
  INVXLTH U11 ( .A(in[6]), .Y(n19) );
  INVXLTH U12 ( .A(in[4]), .Y(n21) );
  INVXLTH U13 ( .A(in[5]), .Y(n20) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U15 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  INVXLTH U16 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U18 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U20 ( .A(in[2]), .Y(n23) );
  NAND2BXLTH U21 ( .AN(in[0]), .B(n17), .Y(out[0]) );
endmodule


module tc_sm_188 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n27, n28, n29, n30, n31, n32, n34, n35,
         n36, n37, n38, n39, n41;

  OA21XLTH U3 ( .A0(in[6]), .A1(n37), .B0(n7), .Y(n27) );
  NAND2XLTH U4 ( .A(n27), .B(n8), .Y(out[3]) );
  CLKINVX12 U5 ( .A(n30), .Y(n8) );
  OR2X2 U6 ( .A(n34), .B(n10), .Y(n28) );
  OR2XLTH U7 ( .A(in[6]), .B(n38), .Y(n29) );
  NAND3XLTH U8 ( .A(n28), .B(n29), .C(n8), .Y(out[2]) );
  OAI221XL U9 ( .A0(n34), .A1(n12), .B0(in[6]), .B1(n39), .C0(n8), .Y(out[1])
         );
  INVXLTH U10 ( .A(in[4]), .Y(n36) );
  INVXLTH U11 ( .A(in[5]), .Y(n35) );
  INVXLTH U12 ( .A(in[6]), .Y(n34) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n37) );
  NOR3X1TH U14 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  AOI21BXLTH U15 ( .A0(n37), .A1(n9), .B0N(in[6]), .Y(n32) );
  INVXLTH U16 ( .A(in[6]), .Y(n31) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U19 ( .A(n38), .B(n11), .Y(n10) );
  NOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U21 ( .A(in[2]), .Y(n38) );
  INVXLTH U22 ( .A(in[1]), .Y(n39) );
  XNOR2XLTH U23 ( .A(in[0]), .B(in[1]), .Y(n12) );
  AOI33X4 U24 ( .A0(n36), .A1(n31), .A2(n35), .B0(n32), .B1(in[4]), .B2(in[5]), 
        .Y(n30) );
  NAND2BXLTH U25 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OA21X4 U18 ( .A0(n9), .A1(n37), .B0(in[6]), .Y(n41) );
  CLKINVX40 U26 ( .A(n41), .Y(n7) );
endmodule


module total_3_test_0 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n61, w5_4_, n5, n6, n7, n8, n43, n44, n45, n50, n51, n52, n53, n54,
         n55, n56, n57;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_191 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_190 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_189 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_188 sm_tc_4 ( .out(in1), .in(in) );
  add_47 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1({a1[6:1], 
        n6}), .in2(b1), .in3(c1), .in(in1) );
  tc_sm_191 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_190 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_189 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_188 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n53), .CK(clk), .RN(n7), 
        .Q(up2[0]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n53), .CK(clk), .RN(n8), 
        .Q(up1[2]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n57), .CK(clk), .RN(n7), .Q(
        h) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n56), .CK(clk), .RN(n7), 
        .Q(up3[3]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n52), .CK(clk), .RN(n7), 
        .Q(n61) );
  SDFFRQXLTH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n54), .CK(clk), .RN(n7), .Q(
        up1[0]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n51), .CK(clk), .RN(n8), 
        .Q(up2[3]) );
  SDFFRQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n54), .CK(clk), .RN(n7), 
        .Q(up1[4]) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n54), .CK(clk), .RN(n7), 
        .Q(up2[4]) );
  SDFFRQXL up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n56), .CK(clk), .RN(n7), 
        .Q(up1[1]) );
  SDFFRQX2 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n53), .CK(clk), .RN(n7), 
        .Q(up3[2]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n53), .CK(clk), .RN(n7), 
        .Q(up3[0]) );
  SDFFRQX1 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n57), .CK(clk), .RN(n7), 
        .Q(up3[1]) );
  INVXLTH U3 ( .A(n5), .Y(n6) );
  INVX2TH U4 ( .A(a1[0]), .Y(n5) );
  CLKBUFX1TH U5 ( .A(rst), .Y(n8) );
  CLKBUFX4TH U6 ( .A(rst), .Y(n7) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n54), .CK(clk), .RN(n7), 
        .Q(up2[1]) );
  SDFFRX4 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n51), .CK(clk), .RN(n7), 
        .Q(up2[2]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n52), .CK(clk), .RN(n8), 
        .Q(up1[3]) );
  INVXLTH U39 ( .A(test_se), .Y(n43) );
  INVXLTH U40 ( .A(n43), .Y(n44) );
  INVXLTH U41 ( .A(n43), .Y(n45) );
  DLY1X1TH U42 ( .A(n55), .Y(n50) );
  INVXLTH U43 ( .A(n50), .Y(n51) );
  INVXLTH U44 ( .A(n50), .Y(n52) );
  DLY1X1TH U45 ( .A(n44), .Y(n53) );
  DLY1X1TH U46 ( .A(n45), .Y(n54) );
  INVXLTH U47 ( .A(n44), .Y(n55) );
  INVXLTH U48 ( .A(n50), .Y(n56) );
  INVXLTH U49 ( .A(n50), .Y(n57) );
  DLY1X1TH U50 ( .A(n61), .Y(up3[4]) );
endmodule


module sm_tc_187 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n26, n27, n30, n31, n32;

  NOR2X4 U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX2 U3 ( .A(in[4]), .Y(n27) );
  OAI2BB2X4 U4 ( .B0(n31), .B1(n6), .A0N(in[1]), .A1N(n31), .Y(out[1]) );
  AOI31X1 U5 ( .A0(n3), .A1(n32), .A2(n5), .B0(n31), .Y(out[4]) );
  CLKBUFX1TH U6 ( .A(out[4]), .Y(out[6]) );
  XNOR2X1TH U7 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U8 ( .A(n8), .B(n26), .Y(n7) );
  CLKBUFX1TH U9 ( .A(in[0]), .Y(out[0]) );
  OAI22XLTH U10 ( .A0(in[4]), .A1(n26), .B0(n31), .B1(n5), .Y(out[2]) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n26) );
  OAI2BB2XLTH U12 ( .B0(n31), .B1(n32), .A0N(in[3]), .A1N(n31), .Y(out[3]) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  AO21XLTH U16 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKINVX40 U15 ( .A(n27), .Y(n30) );
  CLKINVX40 U17 ( .A(n30), .Y(n31) );
  XOR2X1 U18 ( .A(in[2]), .B(n8), .Y(n5) );
  CLKBUFX40 U19 ( .A(n4), .Y(n32) );
endmodule


module sm_tc_186 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n23, n24, n25, n26, n28, n29, n33, n34, n37,
         n38, n39, n40, n41, n42, n43;

  INVX4 U3 ( .A(n23), .Y(n33) );
  BUFX10 U4 ( .A(in[4]), .Y(n23) );
  CLKBUFX1TH U5 ( .A(out[5]), .Y(out[6]) );
  OR2XLTH U7 ( .A(n23), .B(n34), .Y(n24) );
  OR2XLTH U8 ( .A(n33), .B(n5), .Y(n25) );
  NAND2X2 U9 ( .A(n24), .B(n25), .Y(out[2]) );
  INVX8 U10 ( .A(in[2]), .Y(n34) );
  BUFX2 U11 ( .A(n37), .Y(out[0]) );
  NAND2X1 U14 ( .A(n8), .B(n34), .Y(n7) );
  CLKNAND2X2 U15 ( .A(n26), .B(n42), .Y(n29) );
  INVXLTH U16 ( .A(n34), .Y(n26) );
  BUFX2TH U17 ( .A(out[5]), .Y(out[4]) );
  AOI31X4TH U18 ( .A0(n3), .A1(n4), .A2(n5), .B0(n33), .Y(out[5]) );
  CLKNAND2X2 U19 ( .A(n34), .B(n8), .Y(n28) );
  OAI2BB2X1TH U21 ( .B0(n33), .B1(n6), .A0N(in[1]), .A1N(n33), .Y(out[1]) );
  OAI2BB2X1TH U22 ( .B0(n33), .B1(n4), .A0N(in[3]), .A1N(n33), .Y(out[3]) );
  NOR2BXLTH U23 ( .AN(n6), .B(n37), .Y(n3) );
  CLKBUFX40 U2 ( .A(in[0]), .Y(n37) );
  OR2X8 U6 ( .A(in[1]), .B(n37), .Y(n38) );
  CLKINVX40 U12 ( .A(n38), .Y(n8) );
  DLY1X1TH U13 ( .A(n43), .Y(n39) );
  AND2X8 U20 ( .A(n28), .B(n29), .Y(n40) );
  CLKINVX40 U24 ( .A(n40), .Y(n5) );
  AOI21BX4 U25 ( .A0(n37), .A1(in[1]), .B0N(n42), .Y(n41) );
  CLKINVX40 U26 ( .A(n41), .Y(n6) );
  CLKINVX40 U27 ( .A(n8), .Y(n42) );
  XOR2X1 U28 ( .A(n7), .B(in[3]), .Y(n43) );
  CLKINVX40 U29 ( .A(n39), .Y(n4) );
endmodule


module sm_tc_185 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n29, n30, n31, n32, n33, n34, n38, n39, n42,
         n43, n44, n45;

  BUFX8 U2 ( .A(in[4]), .Y(n34) );
  CLKNAND2X8 U4 ( .A(n8), .B(n39), .Y(n7) );
  XNOR2X1TH U5 ( .A(n39), .B(n8), .Y(n5) );
  BUFX5 U7 ( .A(in[0]), .Y(n29) );
  AOI31X4 U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n38), .Y(out[5]) );
  OAI22X2 U9 ( .A0(n34), .A1(n39), .B0(n38), .B1(n5), .Y(out[2]) );
  OAI2BB2X1 U10 ( .B0(n38), .B1(n6), .A0N(in[1]), .A1N(n38), .Y(out[1]) );
  OAI2BB2X4 U11 ( .B0(n38), .B1(n4), .A0N(in[3]), .A1N(n38), .Y(out[3]) );
  INVX4 U12 ( .A(n34), .Y(n38) );
  CLKNAND2X4 U13 ( .A(n32), .B(n33), .Y(n4) );
  INVXLTH U15 ( .A(in[3]), .Y(n31) );
  CLKBUFX1TH U16 ( .A(out[5]), .Y(out[4]) );
  INVX2 U17 ( .A(in[2]), .Y(n39) );
  NAND2X2TH U18 ( .A(n7), .B(in[3]), .Y(n32) );
  INVXL U19 ( .A(n7), .Y(n30) );
  DLY3X1TH U20 ( .A(out[5]), .Y(out[6]) );
  CLKBUFX2TH U21 ( .A(n29), .Y(out[0]) );
  NOR2BXLTH U22 ( .AN(n6), .B(n29), .Y(n3) );
  AOI21BX4 U3 ( .A0(n29), .A1(in[1]), .B0N(n43), .Y(n42) );
  CLKINVX40 U6 ( .A(n42), .Y(n6) );
  CLKINVX40 U14 ( .A(n8), .Y(n43) );
  NOR2BX8 U23 ( .AN(n44), .B(n29), .Y(n8) );
  CLKINVX40 U24 ( .A(in[1]), .Y(n44) );
  AND2X8 U25 ( .A(n30), .B(n31), .Y(n45) );
  CLKINVX40 U26 ( .A(n45), .Y(n33) );
endmodule


module sm_tc_184 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  OAI2BB2X2TH U2 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  OAI2BB2X2TH U3 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKINVX2TH U4 ( .A(in[4]), .Y(n22) );
  CLKBUFX1TH U5 ( .A(in[0]), .Y(out[0]) );
  CLKINVX1TH U6 ( .A(out[4]), .Y(n18) );
  AOI31X4 U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U8 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX1TH U9 ( .A(n18), .Y(out[5]) );
  NOR2X2TH U10 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n21) );
  OAI22X1TH U12 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  INVXLTH U13 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U14 ( .A(n21), .B(n8), .Y(n5) );
  XNOR2X1TH U15 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U16 ( .A(n8), .B(n21), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_46_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  NAND2X2 U1 ( .A(B[1]), .B(n1), .Y(n4) );
  NAND2X1 U2 ( .A(A[1]), .B(B[1]), .Y(n2) );
  AND2X1TH U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  NAND3X2TH U4 ( .A(n2), .B(n3), .C(n4), .Y(carry[2]) );
  CLKNAND2X2TH U5 ( .A(A[1]), .B(n1), .Y(n3) );
  XOR3X1TH U6 ( .A(A[1]), .B(B[1]), .C(n1), .Y(SUM[1]) );
  CLKXOR2X1TH U7 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_46_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  NAND3X2 U1 ( .A(n2), .B(n3), .C(n4), .Y(carry[2]) );
  XOR2XLTH U2 ( .A(n5), .B(carry[3]), .Y(SUM[3]) );
  NAND2X1 U4 ( .A(carry[3]), .B(A[3]), .Y(n6) );
  NAND2X1TH U5 ( .A(A[1]), .B(n9), .Y(n2) );
  NAND3X2 U6 ( .A(n6), .B(n7), .C(n8), .Y(carry[4]) );
  XOR2X2 U7 ( .A(B[5]), .B(A[5]), .Y(n10) );
  NAND2X2 U8 ( .A(carry[5]), .B(A[5]), .Y(n11) );
  NAND2XLTH U9 ( .A(n9), .B(B[1]), .Y(n4) );
  CLKNAND2X2TH U10 ( .A(A[3]), .B(B[3]), .Y(n8) );
  CLKNAND2X2 U11 ( .A(carry[5]), .B(B[5]), .Y(n12) );
  NAND2X2TH U12 ( .A(carry[3]), .B(B[3]), .Y(n7) );
  XOR2X1TH U13 ( .A(B[3]), .B(A[3]), .Y(n5) );
  CLKXOR2X4 U14 ( .A(n10), .B(carry[5]), .Y(SUM[5]) );
  NAND2XLTH U15 ( .A(A[1]), .B(B[1]), .Y(n3) );
  XNOR2X2TH U17 ( .A(n14), .B(A[1]), .Y(SUM[1]) );
  XNOR2XLTH U18 ( .A(B[1]), .B(n9), .Y(n14) );
  CLKXOR2X1TH U19 ( .A(n16), .B(A[0]), .Y(SUM[0]) );
  NAND3X2 U20 ( .A(n11), .B(n12), .C(n13), .Y(carry[6]) );
  AND2X8 U3 ( .A(A[5]), .B(B[5]), .Y(n15) );
  CLKINVX40 U16 ( .A(n15), .Y(n13) );
  DLY1X1TH U21 ( .A(B[0]), .Y(n16) );
  NAND2X8 U22 ( .A(n16), .B(A[0]), .Y(n17) );
  CLKINVX40 U23 ( .A(n17), .Y(n9) );
endmodule


module add_46_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_46_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X4TH U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  XOR2XLTH U2 ( .A(A[6]), .B(B[6]), .Y(n2) );
  AND2XLTH U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_46_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n2, n3, n4, n5, n8, n9, n10, n11, n12, n13;
  wire   [5:2] carry;

  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_4 ( .A(carry[4]), .B(B[4]), .CI(A[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_1 ( .A(n5), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND2X2 U1 ( .A(n8), .B(n9), .Y(SUM[0]) );
  NAND2X1 U2 ( .A(carry[5]), .B(B[5]), .Y(n3) );
  XNOR2X2TH U3 ( .A(n11), .B(carry[5]), .Y(SUM[5]) );
  CLKNAND2X2 U4 ( .A(B[0]), .B(n13), .Y(n8) );
  INVXLTH U5 ( .A(B[0]), .Y(n12) );
  NAND2XLTH U6 ( .A(carry[5]), .B(A[5]), .Y(n2) );
  XNOR2XLTH U7 ( .A(B[5]), .B(A[5]), .Y(n11) );
  NAND2XLTH U8 ( .A(A[5]), .B(B[5]), .Y(n4) );
  CLKNAND2X2 U9 ( .A(n12), .B(A[0]), .Y(n9) );
  INVXLTH U10 ( .A(A[0]), .Y(n13) );
  AND2XLTH U11 ( .A(B[0]), .B(A[0]), .Y(n5) );
  XOR3X2 U12 ( .A(A[6]), .B(B[6]), .C(n10), .Y(SUM[6]) );
  NAND3X2 U13 ( .A(n2), .B(n3), .C(n4), .Y(n10) );
endmodule


module add_46_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR2X3TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_46 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   n28, temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_,
         temp2_0_, temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_,
         temp1_0_, n18, n19, n20, n21, n22, n23, n24, n25, n27;

  add_46_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n27, temp1_0_}), .B({in2[6:2], n25, in2[0]}), .SUM({n28, 
        out3[5:0]}) );
  add_46_DW01_add_1 add_33 ( .A({temp2_6_, n18, temp2_4_, temp2_3_, temp2_2_, 
        n24, temp2_0_}), .B(in), .SUM(out1) );
  add_46_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n27, temp1_0_}), .B({in3[6:3], n23, in3[1:0]}), .SUM(out2)
         );
  add_46_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n27, n22}), .B({temp2_6_, n20, temp2_4_, temp2_3_, temp2_2_, 
        n24, temp2_0_}), .SUM(out) );
  add_46_DW01_add_4 add_30 ( .A({in2[6:2], n25, in2[0]}), .B({in3[6:3], n23, 
        in3[1:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_46_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2 U1 ( .A(in2[1]), .Y(n25) );
  BUFX3 U2 ( .A(temp2_1_), .Y(n24) );
  INVXLTH U3 ( .A(n18), .Y(n19) );
  BUFX10 U4 ( .A(temp2_5_), .Y(n18) );
  CLKBUFX2 U5 ( .A(in3[2]), .Y(n23) );
  INVXLTH U6 ( .A(n19), .Y(n20) );
  INVXLTH U13 ( .A(temp1_0_), .Y(n21) );
  INVXLTH U14 ( .A(n21), .Y(n22) );
  CLKBUFX40 U15 ( .A(n28), .Y(out3[6]) );
  CLKBUFX40 U16 ( .A(temp1_1_), .Y(n27) );
endmodule


module tc_sm_187 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n28, n29, n30, n31, n32, n33;

  CLKBUFX2TH U3 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U4 ( .A(in[1]), .Y(n33) );
  INVXLTH U5 ( .A(in[2]), .Y(n32) );
  XNOR2XLTH U6 ( .A(n32), .B(n11), .Y(n10) );
  INVXLTH U7 ( .A(in[4]), .Y(n30) );
  INVXLTH U8 ( .A(in[5]), .Y(n29) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n31) );
  NAND2BXLTH U10 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI33X4TH U11 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n29), .B2(
        n30), .Y(n8) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U15 ( .A(in[6]), .Y(n28) );
  OAI21XLTH U16 ( .A0(n9), .A1(n31), .B0(in[6]), .Y(n7) );
  OAI221XLTH U17 ( .A0(n28), .A1(n12), .B0(in[6]), .B1(n33), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U18 ( .A0(n28), .A1(n10), .B0(in[6]), .B1(n32), .C0(n8), .Y(
        out[2]) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n31), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n31), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_186 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n21, n22, n23, n24, n25, n26, n28,
         n29, n30, n31, n32, n33, n35;

  CLKINVX1TH U3 ( .A(in[3]), .Y(n31) );
  CLKBUFX1TH U4 ( .A(in[6]), .Y(out[4]) );
  OA21XLTH U5 ( .A0(in[6]), .A1(n31), .B0(n7), .Y(n21) );
  CLKINVX1 U6 ( .A(in[6]), .Y(n28) );
  NAND3XLTH U7 ( .A(n22), .B(n23), .C(n26), .Y(out[2]) );
  NAND3XLTH U8 ( .A(n24), .B(n25), .C(n26), .Y(out[1]) );
  OAI2BB1X4 U9 ( .A0N(n31), .A1N(n9), .B0(in[6]), .Y(n13) );
  NAND2X1 U10 ( .A(n21), .B(n35), .Y(out[3]) );
  OAI21XL U11 ( .A0(n9), .A1(n31), .B0(in[6]), .Y(n7) );
  OR2X1 U12 ( .A(n28), .B(n10), .Y(n22) );
  OR2XLTH U13 ( .A(in[6]), .B(n32), .Y(n23) );
  OR2XL U14 ( .A(n28), .B(n12), .Y(n24) );
  OR2XLTH U15 ( .A(in[6]), .B(n33), .Y(n25) );
  OAI33X4 U16 ( .A0(n13), .A1(n29), .A2(n30), .B0(in[4]), .B1(in[6]), .B2(
        in[5]), .Y(n8) );
  BUFX10 U17 ( .A(n8), .Y(n26) );
  INVXLTH U18 ( .A(in[4]), .Y(n30) );
  INVXLTH U19 ( .A(in[5]), .Y(n29) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n35), .Y(out[0]) );
  INVXLTH U21 ( .A(in[1]), .Y(n33) );
  XNOR2XLTH U22 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U23 ( .A(n32), .B(n11), .Y(n10) );
  NOR2XLTH U24 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U25 ( .A(in[2]), .Y(n32) );
  NOR3X1TH U26 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX40 U27 ( .A(n26), .Y(n35) );
endmodule


module tc_sm_185 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n22, n23, n24, n25, n27, n28,
         n29;

  CLKINVX1TH U4 ( .A(in[3]), .Y(n23) );
  INVXLTH U5 ( .A(in[6]), .Y(n20) );
  NOR3X1TH U6 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U7 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U9 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U10 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U11 ( .A(in[2]), .Y(n24) );
  OAI21XLTH U12 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVX2 U16 ( .A(in[5]), .Y(n21) );
  OAI221XLTH U17 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U18 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(
        out[2]) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
  INVXL U21 ( .A(in[4]), .Y(n22) );
  AOI33X4 U3 ( .A0(n22), .A1(n28), .A2(n21), .B0(n29), .B1(in[5]), .B2(in[4]), 
        .Y(n27) );
  CLKINVX40 U14 ( .A(n27), .Y(n8) );
  CLKINVX40 U20 ( .A(in[6]), .Y(n28) );
  AOI21BX4 U22 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n29) );
endmodule


module tc_sm_184 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n25, n26, n27,
         n28, n29, n30, n32, n33, n34;

  OR3XLTH U6 ( .A(n21), .B(n22), .C(n23), .Y(out[2]) );
  NAND2BXL U7 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OR2XLTH U8 ( .A(n33), .B(n12), .Y(n19) );
  OR2XLTH U9 ( .A(in[6]), .B(n30), .Y(n20) );
  NAND3XLTH U10 ( .A(n19), .B(n20), .C(n8), .Y(out[1]) );
  NOR2XLTH U11 ( .A(n33), .B(n10), .Y(n21) );
  NOR2XLTH U12 ( .A(in[6]), .B(n29), .Y(n22) );
  INVXLTH U13 ( .A(n8), .Y(n23) );
  XNOR2X1TH U14 ( .A(n29), .B(n11), .Y(n10) );
  INVXLTH U15 ( .A(in[6]), .Y(n25) );
  CLKINVX1TH U16 ( .A(in[3]), .Y(n28) );
  NOR3X1TH U17 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U18 ( .A(in[1]), .Y(n30) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U21 ( .A(in[2]), .Y(n29) );
  OAI21XLTH U22 ( .A0(n9), .A1(n28), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U23 ( .A(in[6]), .Y(out[4]) );
  INVX2 U24 ( .A(in[5]), .Y(n26) );
  INVXL U26 ( .A(in[4]), .Y(n27) );
  AOI33X4 U3 ( .A0(n27), .A1(n33), .A2(n26), .B0(n34), .B1(in[5]), .B2(in[4]), 
        .Y(n32) );
  CLKINVX40 U4 ( .A(n32), .Y(n8) );
  CLKINVX40 U5 ( .A(in[6]), .Y(n33) );
  AOI21BX4 U25 ( .A0(n28), .A1(n9), .B0N(in[6]), .Y(n34) );
  OAI2B11X4 U27 ( .A1N(n25), .A0(n28), .B0(n7), .C0(n8), .Y(out[3]) );
endmodule


module total_3_test_1 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n57, n58, w5_4_, n6, n7, n42, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_187 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_186 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_185 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_184 sm_tc_4 ( .out(in1), .in(in) );
  add_46 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_187 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in({n46, w55[5:0]}) );
  tc_sm_186 tc_sm_2 ( .out(w6), .in({n45, w66[5:0]}) );
  tc_sm_185 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_184 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up2[4]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n48), .CK(clk), .RN(n7), .Q(
        h) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n53), .CK(clk), .RN(n7), 
        .Q(n58) );
  SDFFRQXLTH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up1[4]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up3[0]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up2[0]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(n57) );
  SDFFRQXL up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up3[2]) );
  SDFFRQX2 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up1[1]) );
  SDFFRQX2 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n51), .CK(clk), .RN(n7), 
        .Q(up1[2]) );
  SDFFRQX2 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n53), .CK(clk), .RN(n6), 
        .Q(up2[1]) );
  SDFFRQX2 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n54), .CK(clk), .RN(n6), 
        .Q(up2[2]) );
  SDFFRQXL up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up2[3]) );
  SDFFRQX2 up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up3[4]) );
  SDFFRQX2 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up3[1]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n7) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n6) );
  SDFFRX4 up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n54), .CK(clk), .RN(n6), .Q(
        up1[0]) );
  DLY1X1TH U37 ( .A(test_se), .Y(n42) );
  CLKBUFX40 U38 ( .A(w66[6]), .Y(n45) );
  CLKBUFX40 U39 ( .A(w55[6]), .Y(n46) );
  DLY1X1TH U40 ( .A(n52), .Y(n47) );
  INVXLTH U41 ( .A(n47), .Y(n48) );
  INVXLTH U42 ( .A(n47), .Y(n49) );
  DLY1X1TH U43 ( .A(n42), .Y(n50) );
  DLY1X1TH U44 ( .A(n42), .Y(n51) );
  INVXLTH U45 ( .A(n42), .Y(n52) );
  INVXLTH U46 ( .A(n47), .Y(n53) );
  INVXLTH U47 ( .A(n47), .Y(n54) );
  DLY1X1TH U48 ( .A(n57), .Y(up1[3]) );
  DLY1X1TH U49 ( .A(n58), .Y(up3[3]) );
endmodule


module sm_tc_183 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n21, n22;

  INVX2TH U2 ( .A(in[2]), .Y(n22) );
  INVX2 U3 ( .A(in[4]), .Y(n21) );
  BUFX2 U4 ( .A(in[0]), .Y(out[0]) );
  AO21X2 U5 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X4 U6 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKBUFX1TH U7 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX1TH U8 ( .A(out[4]), .Y(out[5]) );
  AOI31X2TH U9 ( .A0(n3), .A1(n4), .A2(n5), .B0(n21), .Y(out[4]) );
  OAI2BB2X4 U10 ( .B0(n21), .B1(n6), .A0N(in[1]), .A1N(n21), .Y(out[1]) );
  XNOR2X2TH U11 ( .A(n22), .B(n8), .Y(n5) );
  XNOR2X4TH U12 ( .A(in[3]), .B(n7), .Y(n4) );
  NAND2XLTH U13 ( .A(n8), .B(n22), .Y(n7) );
  OAI22X1 U14 ( .A0(in[4]), .A1(n22), .B0(n21), .B1(n5), .Y(out[2]) );
  OAI2BB2XLTH U15 ( .B0(n21), .B1(n4), .A0N(in[3]), .A1N(n21), .Y(out[3]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
endmodule


module sm_tc_182 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n23, n24, n25, n27, n30, n31;

  NOR2XLTH U2 ( .A(in[4]), .B(n31), .Y(n23) );
  NOR2X2 U3 ( .A(n30), .B(n5), .Y(n24) );
  OR2X2 U4 ( .A(n23), .B(n24), .Y(out[2]) );
  INVX2 U5 ( .A(in[2]), .Y(n31) );
  INVX2 U6 ( .A(in[4]), .Y(n30) );
  AND2XL U7 ( .A(in[0]), .B(in[1]), .Y(n25) );
  OR2XL U8 ( .A(n25), .B(n8), .Y(n6) );
  OAI2BB2X2 U9 ( .B0(n30), .B1(n6), .A0N(in[1]), .A1N(n30), .Y(out[1]) );
  XNOR2X1TH U10 ( .A(n7), .B(in[3]), .Y(n4) );
  NOR2X6 U11 ( .A(in[1]), .B(in[0]), .Y(n8) );
  AOI31X2TH U12 ( .A0(n3), .A1(n4), .A2(n5), .B0(n30), .Y(out[4]) );
  CLKBUFX1TH U13 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U14 ( .A(n27), .Y(out[6]) );
  NAND2XLTH U15 ( .A(n8), .B(n31), .Y(n7) );
  INVXLTH U16 ( .A(out[4]), .Y(n27) );
  INVXLTH U17 ( .A(n27), .Y(out[5]) );
  NOR2BXLTH U18 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2BB2X1TH U19 ( .B0(n30), .B1(n4), .A0N(in[3]), .A1N(n30), .Y(out[3]) );
  XNOR2X1TH U20 ( .A(n31), .B(n8), .Y(n5) );
endmodule


module sm_tc_181 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n24, n25, n29, n30, n33, n34;

  BUFX20 U2 ( .A(in[4]), .Y(n25) );
  OAI22X2 U3 ( .A0(n25), .A1(n29), .B0(n30), .B1(n5), .Y(out[2]) );
  INVX2 U4 ( .A(n25), .Y(n30) );
  BUFX10 U5 ( .A(in[0]), .Y(out[0]) );
  AOI31X2TH U6 ( .A0(n3), .A1(n24), .A2(n5), .B0(n30), .Y(out[4]) );
  OAI2BB2X4 U8 ( .B0(n30), .B1(n6), .A0N(in[1]), .A1N(n30), .Y(out[1]) );
  NOR2X8 U9 ( .A(in[1]), .B(out[0]), .Y(n8) );
  BUFX10 U10 ( .A(n4), .Y(n24) );
  XNOR2X4 U11 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X1TH U12 ( .B0(n30), .B1(n24), .A0N(in[3]), .A1N(n30), .Y(out[3]) );
  XNOR2X1TH U13 ( .A(n29), .B(n8), .Y(n5) );
  NOR2BXLTH U14 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[6]) );
  INVX2 U18 ( .A(in[2]), .Y(n29) );
  AOI21X8 U7 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n33) );
  CLKINVX40 U17 ( .A(n33), .Y(n6) );
  AND2X8 U19 ( .A(n8), .B(n29), .Y(n34) );
  CLKINVX40 U20 ( .A(n34), .Y(n7) );
endmodule


module sm_tc_180 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  NOR2X3TH U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX2TH U3 ( .A(in[4]), .Y(n22) );
  OAI2BB2X1TH U4 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U5 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1TH U6 ( .A(n7), .B(in[3]), .Y(n4) );
  AOI31X2TH U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  OAI2BB2X1TH U8 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  XNOR2X1TH U9 ( .A(n21), .B(n8), .Y(n5) );
  CLKINVX1TH U10 ( .A(in[2]), .Y(n21) );
  NAND2XLTH U11 ( .A(n8), .B(n21), .Y(n7) );
  NOR2BXLTH U12 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U13 ( .A(out[4]), .Y(n18) );
  INVXLTH U14 ( .A(n18), .Y(out[5]) );
  OAI22X1TH U15 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  INVXLTH U16 ( .A(n18), .Y(out[6]) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_45_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  NAND2XLTH U1 ( .A(A[1]), .B(B[1]), .Y(n3) );
  NAND2X1TH U2 ( .A(B[1]), .B(n1), .Y(n5) );
  NAND2X1TH U3 ( .A(A[1]), .B(n1), .Y(n4) );
  NAND3X2TH U4 ( .A(n3), .B(n4), .C(n5), .Y(carry[2]) );
  CLKXOR2X1TH U5 ( .A(n2), .B(A[1]), .Y(SUM[1]) );
  XOR2XLTH U6 ( .A(n1), .B(B[1]), .Y(n2) );
  CLKXOR2X1TH U7 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1TH U8 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_45_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_45_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_45_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_45_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR2X1 U1 ( .A(B[6]), .B(A[6]), .Y(n2) );
  XOR2X1 U2 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_45_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2TH U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2X2 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_45 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n20, n21, n22, n23, n24, n25, n26, n27;

  add_45_DW01_add_0 add_34 ( .A({temp1_6_, n26, n27, n20, temp1_2_, temp1_1_, 
        temp1_0_}), .B({in2[6:2], n25, in2[0]}), .SUM(out3) );
  add_45_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, n23, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .B({in[6:3], n21, in[1:0]}), .SUM(out1) );
  add_45_DW01_add_2 add_32 ( .A({temp1_6_, n26, n27, n20, temp1_2_, temp1_1_, 
        temp1_0_}), .B({in3[6:2], n24, in3[0]}), .SUM(out2) );
  add_45_DW01_add_3 add_31 ( .A({temp1_6_, n26, n27, n20, temp1_2_, temp1_1_, 
        n22}), .B({temp2_6_, temp2_5_, n23, temp2_3_, temp2_2_, temp2_1_, 
        temp2_0_}), .SUM(out) );
  add_45_DW01_add_4 add_30 ( .A({in2[6:2], n25, in2[0]}), .B({in3[6:2], n24, 
        in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_45_DW01_add_5 add_29 ( .A({in[6:3], n21, in[1:0]}), .B(in1), .SUM({
        temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_})
         );
  BUFX2 U1 ( .A(temp1_3_), .Y(n20) );
  BUFX2TH U2 ( .A(temp2_4_), .Y(n23) );
  CLKBUFX3 U3 ( .A(in3[1]), .Y(n24) );
  BUFX3 U4 ( .A(in2[1]), .Y(n25) );
  BUFX2 U5 ( .A(in[2]), .Y(n21) );
  BUFX2 U6 ( .A(temp1_0_), .Y(n22) );
  CLKBUFX40 U13 ( .A(temp1_5_), .Y(n26) );
  CLKBUFX40 U14 ( .A(temp1_4_), .Y(n27) );
endmodule


module tc_sm_183 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U10 ( .A(in[4]), .Y(n28) );
  INVXLTH U11 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_182 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n21, n22, n23, n26, n27, n28, n29, n31,
         n32;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OR3X2 U3 ( .A(n21), .B(n22), .C(n23), .Y(out[2]) );
  INVX8 U4 ( .A(n6), .Y(n23) );
  OAI211XL U5 ( .A0(in[6]), .A1(n27), .B0(n5), .C0(n6), .Y(out[3]) );
  NOR2XLTH U6 ( .A(n26), .B(n8), .Y(n21) );
  OAI221X1TH U8 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n29), .C0(n6), .Y(out[1]) );
  INVX4 U9 ( .A(in[6]), .Y(n26) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  NOR2XLTH U12 ( .A(in[6]), .B(n28), .Y(n22) );
  OAI21XLTH U14 ( .A0(n7), .A1(n27), .B0(in[6]), .Y(n5) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  XOR2XLTH U16 ( .A(in[0]), .B(n29), .Y(n10) );
  INVXLTH U17 ( .A(in[3]), .Y(n27) );
  INVXLTH U18 ( .A(in[1]), .Y(n29) );
  INVXLTH U19 ( .A(in[2]), .Y(n28) );
  XOR2XLTH U20 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n9) );
  NAND2BXLTH U22 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  AO21X4 U11 ( .A0(in[6]), .A1(n11), .B0(n32), .Y(n31) );
  CLKINVX40 U13 ( .A(n31), .Y(n6) );
  AOI2BB1X4 U23 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n32) );
endmodule


module tc_sm_181 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n26, n27,
         n28;

  OAI221XL U3 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2])
         );
  OAI221XL U4 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1])
         );
  OAI211XLTH U5 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  INVXLTH U8 ( .A(in[6]), .Y(n19) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n22) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U11 ( .A(in[4]), .Y(n21) );
  INVXLTH U12 ( .A(in[5]), .Y(n20) );
  NAND2BXLTH U13 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  XNOR2XLTH U14 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[2]), .Y(n23) );
  INVXLTH U17 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U19 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U20 ( .A(in[6]), .Y(out[4]) );
  AOI33X4 U6 ( .A0(n21), .A1(n27), .A2(n20), .B0(n28), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U7 ( .A(n26), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n27) );
  AOI21BX4 U22 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n28) );
endmodule


module tc_sm_180 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n21, n22, n24, n25, n26, n27;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  AND2X2 U3 ( .A(n22), .B(n21), .Y(n6) );
  INVXL U4 ( .A(in[6]), .Y(n24) );
  OAI221XL U5 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n27), .C0(n6), .Y(out[1])
         );
  OAI21BXL U6 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n21) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  OAI221XLTH U9 ( .A0(n24), .A1(n8), .B0(in[6]), .B1(n26), .C0(n6), .Y(out[2])
         );
  OAI211XLTH U10 ( .A0(in[6]), .A1(n25), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI21XLTH U11 ( .A0(n7), .A1(n25), .B0(in[6]), .Y(n5) );
  INVXLTH U12 ( .A(in[3]), .Y(n25) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  NAND2X1 U15 ( .A(in[6]), .B(n11), .Y(n22) );
  INVXLTH U16 ( .A(in[2]), .Y(n26) );
  XOR2XLTH U17 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n9) );
  XOR2XLTH U19 ( .A(in[0]), .B(n27), .Y(n10) );
  INVXLTH U20 ( .A(in[1]), .Y(n27) );
endmodule


module total_3_test_2 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n4, n5, n6, n7, n8, n9, n44, n51, n52, n53, n54, n55, n56, n57,
         n58;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_183 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_182 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_181 sm_tc_3 ( .out(c1), .in({c[4:2], n6, c[0]}) );
  sm_tc_180 sm_tc_4 ( .out(in1), .in(in) );
  add_45 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1({a1[6:1], 
        n5}), .in2(b1), .in3(c1), .in(in1) );
  tc_sm_183 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_182 tc_sm_2 ( .out(w6), .in({n7, w66[5:0]}) );
  tc_sm_181 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_180 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n55), .CK(clk), .RN(n9), .Q(
        h) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n54), .CK(clk), .RN(n8), .Q(
        up1[0]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n58), .CK(clk), .RN(n8), 
        .Q(up3[0]) );
  SDFFRQXLTH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n53), .CK(clk), .RN(n8), 
        .Q(up2[1]) );
  SDFFRQX1TH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n54), .CK(clk), .RN(n8), 
        .Q(up2[2]) );
  SDFFRQX1TH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n52), .CK(clk), .RN(n9), 
        .Q(up1[2]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n55), .CK(clk), .RN(n8), 
        .Q(up2[4]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n55), .CK(clk), .RN(n8), 
        .Q(up2[0]) );
  SDFFRQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n57), .CK(clk), .RN(n8), 
        .Q(up1[4]) );
  SDFFRQX2 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n58), .CK(clk), .RN(n8), 
        .Q(up3[1]) );
  SDFFRQX1TH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n53), .CK(clk), .RN(n8), 
        .Q(up2[3]) );
  SDFFRQX4 up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n57), .CK(clk), .RN(n9), 
        .Q(up3[4]) );
  BUFX14 U3 ( .A(w66[6]), .Y(n7) );
  CLKBUFX4 U4 ( .A(c[1]), .Y(n6) );
  INVX6 U5 ( .A(a1[0]), .Y(n4) );
  CLKINVX12 U6 ( .A(n4), .Y(n5) );
  CLKBUFX1TH U7 ( .A(rst), .Y(n9) );
  CLKBUFX4TH U8 ( .A(rst), .Y(n8) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n54), .CK(clk), .RN(n8), 
        .Q(up1[1]) );
  SDFFRHQX8 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n54), .CK(clk), .RN(n8), 
        .Q(up3[2]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n52), .CK(clk), .RN(n8), 
        .Q(up1[3]) );
  SDFFRHQX8 up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n55), .CK(clk), .RN(n8), 
        .Q(up3[3]) );
  DLY1X1TH U41 ( .A(test_se), .Y(n44) );
  DLY1X1TH U42 ( .A(n56), .Y(n51) );
  INVXLTH U43 ( .A(n51), .Y(n52) );
  INVXLTH U44 ( .A(n51), .Y(n53) );
  DLY1X1TH U45 ( .A(n44), .Y(n54) );
  DLY1X1TH U46 ( .A(n44), .Y(n55) );
  INVXLTH U47 ( .A(n44), .Y(n56) );
  INVXLTH U48 ( .A(n51), .Y(n57) );
  INVXLTH U49 ( .A(n51), .Y(n58) );
endmodule


module sm_tc_179 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n21, n25, n26;

  OAI22XL U2 ( .A0(n21), .A1(n25), .B0(n26), .B1(n5), .Y(out[2]) );
  XNOR2X2TH U3 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X4 U4 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n26), .Y(out[1]) );
  AO21X4 U5 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  BUFX3 U6 ( .A(in[0]), .Y(out[0]) );
  NOR2X6 U7 ( .A(in[1]), .B(in[0]), .Y(n8) );
  NAND2XL U8 ( .A(n8), .B(n25), .Y(n7) );
  BUFX6 U9 ( .A(in[4]), .Y(n21) );
  INVX4TH U10 ( .A(n21), .Y(n26) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  CLKINVX1TH U12 ( .A(in[2]), .Y(n25) );
  OAI2BB2XLTH U13 ( .B0(n4), .B1(n26), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  AOI31X2TH U14 ( .A0(n3), .A1(n4), .A2(n5), .B0(n26), .Y(out[4]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  XNOR2X1TH U17 ( .A(n25), .B(n8), .Y(n5) );
endmodule


module sm_tc_178 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n27, n28, n31;

  AO21X2 U2 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X6 U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X1 U4 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI22XL U5 ( .A0(in[4]), .A1(n31), .B0(n28), .B1(n5), .Y(out[2]) );
  XNOR2X2 U6 ( .A(n31), .B(n8), .Y(n5) );
  OAI2BB2X2 U7 ( .B0(n28), .B1(n6), .A0N(in[1]), .A1N(n28), .Y(out[1]) );
  NOR2BX2TH U8 ( .AN(n6), .B(in[0]), .Y(n3) );
  AOI31X2TH U9 ( .A0(n3), .A1(n4), .A2(n5), .B0(n28), .Y(out[4]) );
  CLKBUFX1TH U10 ( .A(out[4]), .Y(out[6]) );
  CLKNAND2X2 U11 ( .A(n8), .B(n31), .Y(n7) );
  INVX2TH U12 ( .A(in[4]), .Y(n28) );
  CLKBUFX1TH U13 ( .A(in[0]), .Y(out[0]) );
  CLKINVX1TH U14 ( .A(in[2]), .Y(n27) );
  OAI2BB2X1TH U15 ( .B0(n28), .B1(n4), .A0N(in[3]), .A1N(n28), .Y(out[3]) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX40 U17 ( .A(n27), .Y(n31) );
endmodule


module sm_tc_177 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n28, n32, n33, n36, n37, n38, n39;

  XNOR2X1TH U2 ( .A(n32), .B(n8), .Y(n5) );
  INVX2 U3 ( .A(in[2]), .Y(n32) );
  BUFX2 U5 ( .A(in[4]), .Y(n28) );
  OAI2BB2XL U6 ( .B0(n39), .B1(n4), .A0N(in[3]), .A1N(n39), .Y(out[3]) );
  AOI31X2 U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n39), .Y(out[4]) );
  XNOR2X4 U8 ( .A(n7), .B(in[3]), .Y(n4) );
  NOR2X4 U9 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX2TH U10 ( .A(n28), .Y(n33) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X2TH U12 ( .B0(n39), .B1(n6), .A0N(in[1]), .A1N(n39), .Y(out[1]) );
  BUFX2TH U13 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  AND2X8 U4 ( .A(n8), .B(n32), .Y(n36) );
  CLKINVX40 U16 ( .A(n36), .Y(n7) );
  AOI21X8 U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n37) );
  CLKINVX40 U18 ( .A(n37), .Y(n6) );
  CLKINVX40 U19 ( .A(n33), .Y(n38) );
  CLKINVX40 U20 ( .A(n38), .Y(n39) );
  OAI2BB2X2 U21 ( .B0(n39), .B1(n5), .A0N(n39), .A1N(in[2]), .Y(out[2]) );
endmodule


module sm_tc_176 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n20, n21;

  OAI2BB2X2 U2 ( .B0(n21), .B1(n6), .A0N(in[1]), .A1N(n21), .Y(out[1]) );
  NOR2X2 U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKBUFX1TH U4 ( .A(in[0]), .Y(out[0]) );
  OAI22X1TH U5 ( .A0(in[4]), .A1(n20), .B0(n21), .B1(n5), .Y(out[2]) );
  CLKBUFX1TH U6 ( .A(out[4]), .Y(out[6]) );
  CLKINVX2TH U7 ( .A(in[4]), .Y(n21) );
  CLKINVX1TH U8 ( .A(in[2]), .Y(n20) );
  OAI2BB2X1TH U9 ( .B0(n21), .B1(n4), .A0N(in[3]), .A1N(n21), .Y(out[3]) );
  AOI31X2TH U10 ( .A0(n3), .A1(n4), .A2(n5), .B0(n21), .Y(out[4]) );
  NOR2BXLTH U11 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[5]) );
  XNOR2X1TH U13 ( .A(n20), .B(n8), .Y(n5) );
  XNOR2X1TH U14 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U15 ( .A(n8), .B(n20), .Y(n7) );
  AO21XLTH U16 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_44_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_44_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHX4TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_44_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_44_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_44_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3XL U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(carry[5]), .CI(B[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_44_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n7, n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(n7) );
  ADDFX1TH U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X2 U1 ( .A(n1), .B(A[1]), .Y(n2) );
  CLKXOR2X4 U2 ( .A(n2), .B(B[1]), .Y(SUM[1]) );
  NAND2X4 U3 ( .A(B[1]), .B(A[1]), .Y(n3) );
  NAND2X4 U4 ( .A(B[1]), .B(n1), .Y(n4) );
  NAND2X1 U5 ( .A(A[1]), .B(n1), .Y(n5) );
  NAND3X2 U6 ( .A(n3), .B(n4), .C(n5), .Y(carry[2]) );
  AND2X2 U7 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X2TH U8 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  CLKBUFX40 U9 ( .A(n7), .Y(SUM[5]) );
endmodule


module add_44 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   n25, temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_,
         temp2_0_, temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_,
         temp1_0_, n18, n19, n20, n22, n23, n24;

  add_44_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, n19, n23, temp1_2_, 
        temp1_1_, n22}), .B({in2[6:3], n18, in2[1:0]}), .SUM(out3) );
  add_44_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, n20}), .B(in), .SUM(out1) );
  add_44_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, n19, n23, temp1_2_, 
        temp1_1_, n22}), .B(in3), .SUM({n25, out2[5:0]}) );
  add_44_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, n19, n23, temp1_2_, 
        temp1_1_, n22}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, n20}), .SUM(out) );
  add_44_DW01_add_4 add_30 ( .A({in2[6:3], n24, in2[1:0]}), .B(in3), .SUM({
        temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_})
         );
  add_44_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX1TH U1 ( .A(n24), .Y(n18) );
  CLKBUFX40 U2 ( .A(temp1_4_), .Y(n19) );
  CLKBUFX40 U3 ( .A(temp2_0_), .Y(n20) );
  CLKBUFX40 U4 ( .A(n25), .Y(out2[6]) );
  CLKBUFX40 U5 ( .A(temp1_0_), .Y(n22) );
  CLKBUFX40 U6 ( .A(temp1_3_), .Y(n23) );
  CLKBUFX40 U13 ( .A(in2[2]), .Y(n24) );
endmodule


module tc_sm_179 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n25, n27, n28, n29, n30, n31, n32;

  CLKBUFX2TH U3 ( .A(in[6]), .Y(n25) );
  NOR3X1TH U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U5 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U6 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U7 ( .A(in[2]), .Y(n31) );
  XNOR2XLTH U8 ( .A(n31), .B(n11), .Y(n10) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(n25), .A2(in[5]), .B0(n13), .B1(n28), .B2(
        n29), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n29) );
  INVXLTH U12 ( .A(in[5]), .Y(n28) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n30) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U16 ( .A(n25), .Y(n27) );
  OAI21XLTH U17 ( .A0(n9), .A1(n30), .B0(n25), .Y(n7) );
  OAI221XLTH U18 ( .A0(n27), .A1(n12), .B0(n25), .B1(n32), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U19 ( .A0(n27), .A1(n10), .B0(n25), .B1(n31), .C0(n8), .Y(out[2])
         );
  OAI211XLTH U20 ( .A0(n25), .A1(n30), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U21 ( .A0N(n30), .A1N(n9), .B0(n25), .Y(n13) );
endmodule


module tc_sm_178 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n21, n23, n24, n25, n26, n27,
         n28, n30;

  CLKINVX12 U3 ( .A(n19), .Y(n8) );
  OAI221XL U4 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n27), .C0(n8), .Y(out[2])
         );
  OAI221XL U6 ( .A0(n23), .A1(n12), .B0(in[6]), .B1(n28), .C0(n8), .Y(out[1])
         );
  AOI21BX2 U7 ( .A0(n26), .A1(n9), .B0N(in[6]), .Y(n21) );
  CLKINVX1TH U8 ( .A(in[6]), .Y(n20) );
  OAI21XLTH U9 ( .A0(n9), .A1(n26), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U10 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U11 ( .A(in[5]), .Y(n24) );
  INVXLTH U12 ( .A(in[4]), .Y(n25) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n26) );
  NOR3X1TH U14 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U15 ( .A(n27), .B(n11), .Y(n10) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  AOI33X4 U17 ( .A0(n25), .A1(n20), .A2(n24), .B0(n21), .B1(in[5]), .B2(in[4]), 
        .Y(n19) );
  INVXLTH U18 ( .A(in[1]), .Y(n28) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U21 ( .A(in[2]), .Y(n27) );
  INVXL U22 ( .A(in[6]), .Y(n23) );
  OAI2B11X4 U5 ( .A1N(n30), .A0(n26), .B0(n7), .C0(n8), .Y(out[3]) );
  CLKINVX40 U23 ( .A(in[6]), .Y(n30) );
endmodule


module tc_sm_177 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n18, n19, n20, n21, n22, n25, n26, n27,
         n28, n29, n30, n32, n33, n34;

  NAND3XLTH U4 ( .A(n18), .B(n19), .C(n8), .Y(out[1]) );
  OR3XLTH U5 ( .A(n20), .B(n21), .C(n22), .Y(out[2]) );
  OAI211XL U6 ( .A0(in[6]), .A1(n28), .B0(n7), .C0(n8), .Y(out[3]) );
  OR2X2TH U8 ( .A(n25), .B(n12), .Y(n18) );
  OR2XLTH U9 ( .A(in[6]), .B(n30), .Y(n19) );
  NOR2X1TH U10 ( .A(n25), .B(n10), .Y(n20) );
  NOR2XLTH U11 ( .A(in[6]), .B(n29), .Y(n21) );
  INVXL U12 ( .A(n8), .Y(n22) );
  INVXL U13 ( .A(in[6]), .Y(n25) );
  CLKINVX1TH U14 ( .A(in[3]), .Y(n28) );
  NOR3X1TH U15 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U16 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U18 ( .A(in[1]), .Y(n30) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U20 ( .A(n29), .B(n11), .Y(n10) );
  NOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U22 ( .A(in[2]), .Y(n29) );
  OAI21XLTH U23 ( .A0(n9), .A1(n28), .B0(in[6]), .Y(n7) );
  INVX2 U24 ( .A(in[5]), .Y(n26) );
  INVXL U26 ( .A(in[4]), .Y(n27) );
  AOI33X4 U3 ( .A0(n27), .A1(n33), .A2(n26), .B0(n34), .B1(in[5]), .B2(in[4]), 
        .Y(n32) );
  CLKINVX40 U7 ( .A(n32), .Y(n8) );
  CLKINVX40 U25 ( .A(in[6]), .Y(n33) );
  AOI21BX4 U27 ( .A0(n28), .A1(n9), .B0N(in[6]), .Y(n34) );
endmodule


module tc_sm_176 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n19, n20, n21, n22, n23, n25,
         n26, n27, n28, n29, n30, n32, n33;

  OAI2BB1X1 U3 ( .A0N(n28), .A1N(n9), .B0(in[6]), .Y(n13) );
  BUFX6 U5 ( .A(n8), .Y(n23) );
  NAND2XLTH U6 ( .A(n18), .B(n23), .Y(out[3]) );
  OA21XL U8 ( .A0(in[6]), .A1(n28), .B0(n7), .Y(n18) );
  INVX2TH U9 ( .A(in[3]), .Y(n28) );
  OR2X2TH U10 ( .A(n25), .B(n12), .Y(n19) );
  OR2XLTH U11 ( .A(in[6]), .B(n30), .Y(n20) );
  OR2X1 U12 ( .A(n25), .B(n10), .Y(n21) );
  OR2XLTH U13 ( .A(in[6]), .B(n29), .Y(n22) );
  INVXL U14 ( .A(in[6]), .Y(n25) );
  NOR3X1TH U15 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U16 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U17 ( .A(in[1]), .Y(n30) );
  XNOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U19 ( .A(n29), .B(n11), .Y(n10) );
  NOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U21 ( .A(in[2]), .Y(n29) );
  OAI21XLTH U22 ( .A0(n9), .A1(n28), .B0(in[6]), .Y(n7) );
  NAND2BXLTH U23 ( .AN(in[0]), .B(n23), .Y(out[0]) );
  OAI33X4 U24 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n26), .B2(
        n27), .Y(n8) );
  INVXL U25 ( .A(in[5]), .Y(n26) );
  INVXL U26 ( .A(in[4]), .Y(n27) );
  AND3X8 U4 ( .A(n21), .B(n22), .C(n23), .Y(n32) );
  CLKINVX40 U7 ( .A(n32), .Y(out[2]) );
  AND3X8 U27 ( .A(n19), .B(n20), .C(n23), .Y(n33) );
  CLKINVX40 U28 ( .A(n33), .Y(out[1]) );
endmodule


module total_3_test_3 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n64, w5_4_, n4, n5, n40, n48, n49, n50, n51, n52, n53, n54, n55;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_179 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_178 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_177 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_176 sm_tc_4 ( .out(in1), .in(in) );
  add_44 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_179 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_178 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_177 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_176 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(n64) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n55), .CK(clk), .RN(n5), .Q(
        h) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up2[3]) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQXLTH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n52), .CK(clk), .RN(n4), .Q(
        up1[0]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  SDFFRQX2 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n52), .CK(clk), .RN(n5), 
        .Q(up1[2]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n5) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n4) );
  SDFFRX4 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n55), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  SDFFRX4 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRX4 up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n54), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRX4 up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up3[3]) );
  SDFFRHQX8 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n54), .CK(clk), .RN(n4), 
        .Q(up1[1]) );
  DLY1X1TH U37 ( .A(test_se), .Y(n40) );
  DLY1X1TH U38 ( .A(n53), .Y(n48) );
  INVXLTH U39 ( .A(n48), .Y(n49) );
  INVXLTH U40 ( .A(n48), .Y(n50) );
  DLY1X1TH U41 ( .A(n40), .Y(n51) );
  DLY1X1TH U42 ( .A(n40), .Y(n52) );
  INVXLTH U43 ( .A(n40), .Y(n53) );
  INVXLTH U44 ( .A(n48), .Y(n54) );
  INVXLTH U45 ( .A(n48), .Y(n55) );
  DLY1X1TH U46 ( .A(n64), .Y(up1[4]) );
endmodule


module sm_tc_175 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n24, n25, n26, n29, n30, n33, n34, n35,
         n36, n37, n38, n39;

  CLKINVX12 U2 ( .A(n22), .Y(out[0]) );
  XNOR2X4 U3 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2X2 U4 ( .A(n8), .B(n29), .Y(n7) );
  NAND2X6 U5 ( .A(n25), .B(n26), .Y(n5) );
  OAI2BB2X4 U6 ( .B0(n38), .B1(n6), .A0N(in[1]), .A1N(n38), .Y(out[1]) );
  NAND2X4 U7 ( .A(in[2]), .B(n24), .Y(n26) );
  OAI22XLTH U9 ( .A0(n37), .A1(n29), .B0(n38), .B1(n5), .Y(out[2]) );
  INVX2 U10 ( .A(in[0]), .Y(n22) );
  INVX4TH U12 ( .A(in[2]), .Y(n29) );
  CLKINVX1TH U13 ( .A(n8), .Y(n24) );
  AOI31X1 U14 ( .A0(n3), .A1(n4), .A2(n5), .B0(n38), .Y(out[4]) );
  INVX3TH U15 ( .A(in[4]), .Y(n30) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2XLTH U17 ( .B0(n38), .B1(n4), .A0N(in[3]), .A1N(n38), .Y(out[3]) );
  CLKBUFX1TH U18 ( .A(out[4]), .Y(out[5]) );
  AO21X2 U19 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OR2X8 U8 ( .A(n34), .B(out[0]), .Y(n33) );
  CLKINVX40 U11 ( .A(n33), .Y(n3) );
  CLKINVX40 U20 ( .A(n6), .Y(n34) );
  NAND2BX8 U21 ( .AN(in[1]), .B(n22), .Y(n35) );
  CLKINVX40 U22 ( .A(n35), .Y(n8) );
  CLKBUFX40 U23 ( .A(n30), .Y(n36) );
  CLKINVX40 U24 ( .A(n36), .Y(n37) );
  CLKINVX40 U25 ( .A(n37), .Y(n38) );
  AND2X8 U26 ( .A(n29), .B(n8), .Y(n39) );
  CLKINVX40 U27 ( .A(n39), .Y(n25) );
endmodule


module sm_tc_174 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n37, n40, n41, n44;

  AOI31X2 U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n40), .Y(out[4]) );
  NAND2X2 U3 ( .A(n34), .B(n35), .Y(n5) );
  OAI2BB2X4TH U4 ( .B0(n40), .B1(n4), .A0N(in[3]), .A1N(n40), .Y(out[3]) );
  INVX6 U5 ( .A(out[4]), .Y(n37) );
  BUFX10 U6 ( .A(in[4]), .Y(n29) );
  CLKNAND2X8 U7 ( .A(n27), .B(n28), .Y(n4) );
  NAND2X4 U8 ( .A(n25), .B(n26), .Y(n28) );
  INVXLTH U9 ( .A(in[3]), .Y(n26) );
  INVXLTH U10 ( .A(n7), .Y(n25) );
  INVX2 U12 ( .A(in[2]), .Y(n41) );
  NAND2X2 U13 ( .A(n7), .B(in[3]), .Y(n27) );
  NAND2X1TH U14 ( .A(n8), .B(n41), .Y(n7) );
  NAND2XL U15 ( .A(n41), .B(n8), .Y(n34) );
  INVXLTH U16 ( .A(n8), .Y(n33) );
  AO21X4 U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  INVX4 U18 ( .A(n29), .Y(n40) );
  CLKBUFX3 U19 ( .A(in[0]), .Y(out[0]) );
  NOR2XL U20 ( .A(n29), .B(n41), .Y(n30) );
  NOR2X8 U21 ( .A(n40), .B(n5), .Y(n31) );
  OR2X8 U22 ( .A(n30), .B(n31), .Y(out[2]) );
  CLKNAND2X4 U23 ( .A(n32), .B(n33), .Y(n35) );
  INVXLTH U24 ( .A(n41), .Y(n32) );
  NOR2BXLTH U25 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U26 ( .A(n37), .Y(out[5]) );
  OAI2BB2X2 U27 ( .B0(n40), .B1(n6), .A0N(in[1]), .A1N(n40), .Y(out[1]) );
  INVXLTH U28 ( .A(n37), .Y(out[6]) );
  OR2X8 U11 ( .A(in[1]), .B(in[0]), .Y(n44) );
  CLKINVX40 U29 ( .A(n44), .Y(n8) );
endmodule


module sm_tc_173 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n23, n24, n28, n29, n32;

  OAI2BB2X4 U2 ( .B0(n28), .B1(n4), .A0N(in[3]), .A1N(n28), .Y(out[3]) );
  BUFX10 U3 ( .A(in[4]), .Y(n24) );
  OAI22X1 U5 ( .A0(n24), .A1(n29), .B0(n28), .B1(n5), .Y(out[2]) );
  AOI31X2 U6 ( .A0(n3), .A1(n4), .A2(n5), .B0(n28), .Y(out[4]) );
  AND2X2 U7 ( .A(out[0]), .B(in[1]), .Y(n23) );
  OR2X2 U8 ( .A(n23), .B(n8), .Y(n6) );
  BUFX5 U9 ( .A(in[0]), .Y(out[0]) );
  NOR2X2 U10 ( .A(in[1]), .B(out[0]), .Y(n8) );
  OAI2BB2X2 U11 ( .B0(n28), .B1(n6), .A0N(in[1]), .A1N(n28), .Y(out[1]) );
  INVX3TH U13 ( .A(n24), .Y(n28) );
  XNOR2X1 U14 ( .A(n29), .B(n8), .Y(n5) );
  INVX1TH U15 ( .A(in[2]), .Y(n29) );
  NOR2BXLTH U16 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U18 ( .A(out[4]), .Y(out[6]) );
  XOR2X1 U4 ( .A(n32), .B(in[3]), .Y(n4) );
  CLKAND2X12 U12 ( .A(n8), .B(n29), .Y(n32) );
endmodule


module sm_tc_172 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  OAI2BB2X2 U2 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  AOI31X4 U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  XNOR2X1TH U4 ( .A(n7), .B(in[3]), .Y(n4) );
  NOR2X2TH U5 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI22X1TH U6 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  OAI2BB2X1TH U7 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U8 ( .A(in[0]), .Y(out[0]) );
  CLKINVX1TH U9 ( .A(in[2]), .Y(n21) );
  CLKINVX2TH U10 ( .A(in[4]), .Y(n22) );
  INVXLTH U11 ( .A(out[4]), .Y(n18) );
  NOR2BXLTH U12 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U13 ( .A(n18), .Y(out[5]) );
  INVXLTH U14 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U15 ( .A(n21), .B(n8), .Y(n5) );
  NAND2XLTH U16 ( .A(n8), .B(n21), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_43_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_43_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [6:2] carry;

  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CLKXOR2X8 U1 ( .A(n6), .B(carry[6]), .Y(SUM[6]) );
  NAND3X4 U3 ( .A(n3), .B(n4), .C(n5), .Y(carry[5]) );
  CLKXOR2X4 U6 ( .A(n2), .B(carry[4]), .Y(SUM[4]) );
  CLKNAND2X2 U7 ( .A(A[4]), .B(B[4]), .Y(n5) );
  CLKXOR2X1TH U8 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X4 U9 ( .A(B[6]), .B(A[6]), .Y(n6) );
  XOR2XLTH U10 ( .A(B[4]), .B(A[4]), .Y(n2) );
  AND2X8 U2 ( .A(carry[4]), .B(B[4]), .Y(n7) );
  CLKINVX40 U4 ( .A(n7), .Y(n4) );
  NAND2X8 U5 ( .A(B[0]), .B(A[0]), .Y(n8) );
  CLKINVX40 U11 ( .A(n8), .Y(n1) );
  AND2X8 U12 ( .A(carry[4]), .B(A[4]), .Y(n9) );
  CLKINVX40 U13 ( .A(n9), .Y(n3) );
endmodule


module add_43_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X8TH U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X4 U3 ( .A(B[6]), .B(A[6]), .Y(n2) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_43_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX4TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_43_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [6:2] carry;

  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n8), .CO(carry[2]), .S(SUM[1]) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR2X1 U1 ( .A(A[3]), .B(B[3]), .Y(n9) );
  CLKXOR2X2 U2 ( .A(n9), .B(carry[3]), .Y(SUM[3]) );
  NAND3X2 U3 ( .A(n5), .B(n6), .C(n7), .Y(carry[4]) );
  NAND2X2 U4 ( .A(n3), .B(n4), .Y(SUM[0]) );
  NAND2XLTH U5 ( .A(A[3]), .B(B[3]), .Y(n7) );
  NAND2XLTH U6 ( .A(carry[3]), .B(A[3]), .Y(n5) );
  NAND2XLTH U7 ( .A(n10), .B(A[0]), .Y(n4) );
  NAND2XLTH U8 ( .A(carry[3]), .B(B[3]), .Y(n6) );
  INVXLTH U9 ( .A(A[0]), .Y(n11) );
  AND2XLTH U11 ( .A(B[0]), .B(A[0]), .Y(n8) );
  INVXLTH U12 ( .A(B[0]), .Y(n10) );
  AND2X8 U10 ( .A(B[0]), .B(n11), .Y(n12) );
  CLKINVX40 U13 ( .A(n12), .Y(n3) );
endmodule


module add_43_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR2XL U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_43 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32;

  add_43_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n32, temp1_2_, 
        temp1_1_, n31}), .B({in2[6:3], n23, n28, in2[0]}), .SUM(out3) );
  add_43_DW01_add_1 add_33 ( .A({n29, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, n22}), .B(in), .SUM(out1) );
  add_43_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n32, temp1_2_, 
        temp1_1_, n31}), .B({n27, in3[5:0]}), .SUM(out2) );
  add_43_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n32, temp1_2_, 
        temp1_1_, n31}), .B({n29, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, n22}), .SUM(out) );
  add_43_DW01_add_4 add_30 ( .A({in2[6:3], n23, n28, in2[0]}), .B({n27, 
        in3[5:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_43_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  INVX2TH U1 ( .A(n21), .Y(n22) );
  INVX2 U2 ( .A(temp2_0_), .Y(n21) );
  INVX2TH U3 ( .A(n24), .Y(n25) );
  INVXLTH U4 ( .A(temp1_0_), .Y(n24) );
  BUFX20 U5 ( .A(in2[2]), .Y(n23) );
  INVXLTH U6 ( .A(n26), .Y(n27) );
  INVXLTH U13 ( .A(in3[6]), .Y(n26) );
  CLKBUFX40 U14 ( .A(in2[1]), .Y(n28) );
  CLKBUFX40 U15 ( .A(temp2_6_), .Y(n29) );
  CLKINVX40 U16 ( .A(n25), .Y(n30) );
  CLKINVX40 U17 ( .A(n30), .Y(n31) );
  CLKBUFX40 U18 ( .A(temp1_3_), .Y(n32) );
endmodule


module tc_sm_175 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U10 ( .A(in[5]), .Y(n27) );
  INVXLTH U11 ( .A(in[4]), .Y(n28) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_174 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n33, n34, n36, n37, n38,
         n39, n41, n42, n43;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  AOI2BB1X2 U3 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  OAI211XL U4 ( .A0(in[6]), .A1(n37), .B0(n5), .C0(n6), .Y(out[3]) );
  OR2XLTH U9 ( .A(n36), .B(n10), .Y(n33) );
  NOR2X1 U11 ( .A(n36), .B(n8), .Y(n30) );
  NOR2XL U12 ( .A(in[6]), .B(n38), .Y(n31) );
  CLKINVX1 U13 ( .A(in[6]), .Y(n36) );
  OAI21XL U14 ( .A0(n7), .A1(n37), .B0(in[6]), .Y(n5) );
  INVXLTH U15 ( .A(in[1]), .Y(n39) );
  NOR3X1TH U16 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  XOR2XLTH U17 ( .A(in[0]), .B(n39), .Y(n10) );
  INVXLTH U18 ( .A(in[3]), .Y(n37) );
  XOR2XLTH U19 ( .A(in[2]), .B(n9), .Y(n8) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  CLKBUFX1TH U21 ( .A(in[6]), .Y(out[4]) );
  OR2XLTH U22 ( .A(in[6]), .B(n39), .Y(n34) );
  INVXLTH U23 ( .A(in[2]), .Y(n38) );
  NOR2XLTH U24 ( .A(in[0]), .B(in[1]), .Y(n9) );
  AND3X8 U5 ( .A(n33), .B(n34), .C(n6), .Y(n41) );
  CLKINVX40 U6 ( .A(n41), .Y(out[1]) );
  NOR3X8 U8 ( .A(n30), .B(n31), .C(n43), .Y(n42) );
  CLKINVX40 U10 ( .A(n42), .Y(out[2]) );
  AO21X4 U25 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n43) );
  CLKINVX40 U26 ( .A(n43), .Y(n6) );
endmodule


module tc_sm_173 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n21, n22, n23, n24, n25, n26, n28, n29,
         n30;

  INVXLTH U4 ( .A(in[5]), .Y(n22) );
  OAI211XLTH U5 ( .A0(in[6]), .A1(n24), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221XLTH U6 ( .A0(n21), .A1(n12), .B0(in[6]), .B1(n26), .C0(n8), .Y(out[1]) );
  OAI221X1TH U7 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[2]) );
  INVX2TH U8 ( .A(in[4]), .Y(n23) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n24) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U11 ( .A(n25), .B(n11), .Y(n10) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U13 ( .A(in[2]), .Y(n25) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U19 ( .A0(n9), .A1(n24), .B0(in[6]), .Y(n7) );
  INVXLTH U20 ( .A(in[6]), .Y(n21) );
  AOI33X4 U3 ( .A0(n23), .A1(n29), .A2(n22), .B0(n30), .B1(in[5]), .B2(in[4]), 
        .Y(n28) );
  CLKINVX40 U18 ( .A(n28), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n29) );
  AOI21BX4 U22 ( .A0(n24), .A1(n9), .B0N(in[6]), .Y(n30) );
endmodule


module tc_sm_172 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n19, n21, n22, n23, n24, n25,
         n26;

  OA21XL U3 ( .A0(in[6]), .A1(n24), .B0(n7), .Y(n18) );
  NAND2XL U4 ( .A(n18), .B(n19), .Y(out[3]) );
  OAI21XL U5 ( .A0(n9), .A1(n24), .B0(in[6]), .Y(n7) );
  OAI33X4 U6 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n22), .B2(n23), .Y(n8) );
  OAI2BB1X4 U7 ( .A0N(n24), .A1N(n9), .B0(in[6]), .Y(n13) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n24) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U10 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U11 ( .A(n25), .B(n11), .Y(n10) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U13 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U15 ( .A(in[6]), .Y(n21) );
  BUFX10 U16 ( .A(n8), .Y(n19) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n19), .Y(out[0]) );
  INVX2 U18 ( .A(in[5]), .Y(n22) );
  OAI221XLTH U19 ( .A0(n21), .A1(n12), .B0(in[6]), .B1(n26), .C0(n19), .Y(
        out[1]) );
  OAI221XLTH U20 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n25), .C0(n19), .Y(
        out[2]) );
  INVXLTH U21 ( .A(in[2]), .Y(n25) );
  INVXL U22 ( .A(in[4]), .Y(n23) );
endmodule


module total_3_test_4 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n4, n5, n40, n45, n46, n47, n48, n49, n50, n51, n52;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_175 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_174 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_173 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_172 sm_tc_4 ( .out(in1), .in(in) );
  add_43 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_175 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_174 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_173 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_172 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n52), .CK(clk), .RN(n4), .Q(
        up1[0]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n46), .CK(clk), .RN(n5), .Q(
        h) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRHQX2TH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  SDFFRHQX2TH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up2[3]) );
  SDFFRQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up1[4]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up3[3]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up1[2]) );
  SDFFRQXL up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  SDFFRQX2 up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  CLKBUFX4TH U3 ( .A(rst), .Y(n4) );
  CLKBUFX1TH U4 ( .A(rst), .Y(n5) );
  SDFFRX4 up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n46), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  INVXLTH U37 ( .A(n50), .Y(n40) );
  DLY1X1TH U38 ( .A(n50), .Y(n45) );
  INVXLTH U39 ( .A(n45), .Y(n46) );
  INVXLTH U40 ( .A(n45), .Y(n47) );
  DLY1X1TH U41 ( .A(n40), .Y(n48) );
  DLY1X1TH U42 ( .A(test_se), .Y(n49) );
  INVXLTH U43 ( .A(test_se), .Y(n50) );
  INVXLTH U44 ( .A(n45), .Y(n51) );
  INVXLTH U45 ( .A(n45), .Y(n52) );
endmodule


module sm_tc_171 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n23, n26;

  INVX2TH U2 ( .A(in[2]), .Y(n23) );
  CLKBUFX1TH U3 ( .A(out[4]), .Y(out[6]) );
  XNOR2X2 U5 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX4 U6 ( .A(in[4]), .Y(n22) );
  AO21X1 U7 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  AOI31X1 U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  OAI2BB2X1 U9 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  OAI2BB2X4TH U10 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  OAI22X2 U12 ( .A0(in[4]), .A1(n23), .B0(n22), .B1(n5), .Y(out[2]) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  NAND2XLTH U15 ( .A(n8), .B(n23), .Y(n7) );
  BUFX2TH U16 ( .A(in[0]), .Y(out[0]) );
  OR2X8 U4 ( .A(in[1]), .B(in[0]), .Y(n26) );
  CLKINVX40 U11 ( .A(n26), .Y(n8) );
  XOR2X1 U17 ( .A(n23), .B(n26), .Y(n5) );
endmodule


module sm_tc_170 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n38, n3, n4, n5, n6, n8, n30, n31, n33, n34, n35, n36;

  OAI22X1 U11 ( .A0(in[4]), .A1(n30), .B0(n35), .B1(n5), .Y(out[2]) );
  CLKBUFX3 U2 ( .A(out[6]), .Y(out[4]) );
  CLKBUFX2TH U3 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X1 U5 ( .B0(n35), .B1(n6), .A0N(in[1]), .A1N(n35), .Y(out[1]) );
  NOR2X4 U6 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI2BB2X1TH U7 ( .B0(n35), .B1(n4), .A0N(in[3]), .A1N(n35), .Y(out[3]) );
  AOI31X2TH U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n35), .Y(n38) );
  INVX2TH U9 ( .A(in[4]), .Y(n31) );
  CLKBUFX1TH U10 ( .A(out[6]), .Y(out[5]) );
  NOR2BXLTH U12 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVX2 U14 ( .A(in[2]), .Y(n30) );
  AO21XLTH U15 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  XNOR2X1TH U16 ( .A(n30), .B(n8), .Y(n5) );
  XOR2X1 U4 ( .A(n33), .B(in[3]), .Y(n4) );
  CLKAND2X12 U13 ( .A(n8), .B(n30), .Y(n33) );
  CLKINVX40 U17 ( .A(n31), .Y(n34) );
  CLKINVX40 U18 ( .A(n34), .Y(n35) );
  CLKINVX40 U19 ( .A(n38), .Y(n36) );
  CLKINVX40 U20 ( .A(n36), .Y(out[6]) );
endmodule


module sm_tc_169 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n26, n27, n29;

  OAI22XL U2 ( .A0(in[4]), .A1(n26), .B0(n27), .B1(n5), .Y(out[2]) );
  AOI31X4 U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n27), .Y(out[6]) );
  XNOR2X1 U4 ( .A(n26), .B(n8), .Y(n5) );
  XNOR2X1TH U6 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKINVX4 U7 ( .A(in[4]), .Y(n27) );
  OAI2BB2X4 U8 ( .B0(n27), .B1(n6), .A0N(in[1]), .A1N(n27), .Y(out[1]) );
  OAI2BB2X2TH U9 ( .B0(n27), .B1(n4), .A0N(in[3]), .A1N(n27), .Y(out[3]) );
  AO21XLTH U10 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2BXLTH U11 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U12 ( .A(out[6]), .Y(out[5]) );
  CLKBUFX1TH U13 ( .A(out[6]), .Y(out[4]) );
  NAND2XLTH U14 ( .A(n8), .B(n26), .Y(n7) );
  BUFX2TH U15 ( .A(in[0]), .Y(out[0]) );
  INVX2 U16 ( .A(in[2]), .Y(n26) );
  OR2X8 U5 ( .A(in[1]), .B(in[0]), .Y(n29) );
  CLKINVX40 U17 ( .A(n29), .Y(n8) );
endmodule


module sm_tc_168 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  NOR2X2 U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  AOI31X2TH U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  OAI22X2TH U4 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  OAI2BB2X1TH U5 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  XNOR2X2TH U6 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX1TH U7 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U8 ( .A(n18), .Y(out[6]) );
  OAI2BB2X2TH U9 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKINVX1TH U10 ( .A(in[2]), .Y(n21) );
  CLKINVX2TH U11 ( .A(in[4]), .Y(n22) );
  INVXLTH U12 ( .A(out[4]), .Y(n18) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U14 ( .A(n18), .Y(out[5]) );
  XNOR2X1TH U15 ( .A(n21), .B(n8), .Y(n5) );
  NAND2XLTH U16 ( .A(n8), .B(n21), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_42_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CLKXOR2X8 U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  XOR2X1TH U2 ( .A(B[6]), .B(A[6]), .Y(n2) );
  AND2XLTH U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_42_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_42_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_42_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_42_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHX2TH U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_42_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n3, n1;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X4TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1 U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(n3) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  CLKBUFX40 U3 ( .A(n3), .Y(SUM[1]) );
endmodule


module add_42 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n27, n29, n30;

  add_42_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n30, 
        temp1_1_, temp1_0_}), .B(in2), .SUM(out3) );
  add_42_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, n29}), .B(in), .SUM(out1) );
  add_42_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n30, 
        temp1_1_, temp1_0_}), .B({in3[6:3], n27, in3[1:0]}), .SUM(out2) );
  add_42_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n30, 
        temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, n29}), .SUM(out) );
  add_42_DW01_add_4 add_30 ( .A(in2), .B({in3[6:3], n27, in3[1:0]}), .SUM({
        temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_})
         );
  add_42_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2 U1 ( .A(in3[2]), .Y(n27) );
  CLKBUFX40 U2 ( .A(temp2_0_), .Y(n29) );
  CLKBUFX40 U3 ( .A(temp1_2_), .Y(n30) );
endmodule


module tc_sm_171 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29, n30;

  CLKBUFX1TH U3 ( .A(in[6]), .Y(out[4]) );
  CLKBUFX2TH U4 ( .A(in[6]), .Y(n24) );
  NOR3X1TH U5 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U6 ( .A(in[1]), .Y(n30) );
  XNOR2XLTH U7 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U8 ( .A(in[2]), .Y(n29) );
  XNOR2XLTH U9 ( .A(n29), .B(n11), .Y(n10) );
  NOR2XLTH U10 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U11 ( .A(n24), .Y(n25) );
  OAI33X4TH U12 ( .A0(in[4]), .A1(n24), .A2(in[5]), .B0(n13), .B1(n26), .B2(
        n27), .Y(n8) );
  INVXLTH U13 ( .A(in[4]), .Y(n27) );
  INVXLTH U14 ( .A(in[5]), .Y(n26) );
  CLKINVX1TH U15 ( .A(in[3]), .Y(n28) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U17 ( .A0(n25), .A1(n12), .B0(n24), .B1(n30), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U18 ( .A0(n25), .A1(n10), .B0(n24), .B1(n29), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U19 ( .A0(n9), .A1(n28), .B0(n24), .Y(n7) );
  OAI211XLTH U20 ( .A0(n24), .A1(n28), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U21 ( .A0N(n28), .A1N(n9), .B0(n24), .Y(n13) );
endmodule


module tc_sm_170 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n31, n32, n33, n34, n36, n37;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OAI211XL U3 ( .A0(n37), .A1(n32), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI221XL U5 ( .A0(n31), .A1(n8), .B0(n37), .B1(n33), .C0(n6), .Y(out[2]) );
  INVXLTH U6 ( .A(in[6]), .Y(n31) );
  OAI221XL U8 ( .A0(n31), .A1(n10), .B0(n37), .B1(n34), .C0(n6), .Y(out[1]) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  NOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI21XLTH U12 ( .A0(n7), .A1(n32), .B0(n37), .Y(n5) );
  CLKBUFX1TH U13 ( .A(n37), .Y(out[4]) );
  XOR2XLTH U14 ( .A(in[0]), .B(n34), .Y(n10) );
  INVXLTH U15 ( .A(in[1]), .Y(n34) );
  INVXLTH U16 ( .A(in[3]), .Y(n32) );
  INVXLTH U17 ( .A(in[2]), .Y(n33) );
  XOR2XLTH U18 ( .A(in[2]), .B(n9), .Y(n8) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  AOI21X8 U4 ( .A0(n37), .A1(n11), .B0(n36), .Y(n6) );
  AOI2BB1X4 U9 ( .A0N(in[5]), .A1N(in[4]), .B0(n37), .Y(n36) );
  CLKBUFX40 U20 ( .A(in[6]), .Y(n37) );
endmodule


module tc_sm_169 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n17, n18, n19, n20, n22, n23, n24, n25,
         n26, n27, n29;

  AOI33X2 U3 ( .A0(n24), .A1(n18), .A2(n23), .B0(n19), .B1(in[5]), .B2(in[4]), 
        .Y(n17) );
  CLKINVX40 U4 ( .A(n29), .Y(n8) );
  CLKINVX40 U5 ( .A(in[6]), .Y(n18) );
  AOI21BX2 U6 ( .A0(n25), .A1(n9), .B0N(in[6]), .Y(n19) );
  OAI221XL U7 ( .A0(n22), .A1(n12), .B0(in[6]), .B1(n27), .C0(n8), .Y(out[1])
         );
  OAI221XL U8 ( .A0(n22), .A1(n10), .B0(in[6]), .B1(n26), .C0(n8), .Y(out[2])
         );
  OA21XLTH U9 ( .A0(in[6]), .A1(n25), .B0(n7), .Y(n20) );
  NAND2XLTH U10 ( .A(n20), .B(n8), .Y(out[3]) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n25) );
  INVXLTH U12 ( .A(in[6]), .Y(n22) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U15 ( .A0(n9), .A1(n25), .B0(in[6]), .Y(n7) );
  XNOR2XLTH U16 ( .A(n26), .B(n11), .Y(n10) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U18 ( .A(in[1]), .Y(n27) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U21 ( .A(in[2]), .Y(n26) );
  INVXL U22 ( .A(in[5]), .Y(n23) );
  INVXL U23 ( .A(in[4]), .Y(n24) );
  CLKBUFX40 U24 ( .A(n17), .Y(n29) );
endmodule


module tc_sm_168 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n18, n19, n21, n22, n23, n24, n25, n26,
         n28, n29, n30;

  OAI211XL U4 ( .A0(in[6]), .A1(n24), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221XL U5 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[2])
         );
  NAND3XL U6 ( .A(n18), .B(n19), .C(n8), .Y(out[1]) );
  OR2XLTH U7 ( .A(n21), .B(n12), .Y(n18) );
  OR2XLTH U8 ( .A(in[6]), .B(n26), .Y(n19) );
  INVXLTH U9 ( .A(in[4]), .Y(n23) );
  INVX1TH U10 ( .A(in[5]), .Y(n22) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n24) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U13 ( .A(n25), .B(n11), .Y(n10) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U16 ( .A0(n9), .A1(n24), .B0(in[6]), .Y(n7) );
  INVXLTH U17 ( .A(in[6]), .Y(n21) );
  INVXLTH U18 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U21 ( .A(in[2]), .Y(n25) );
  AOI33X4 U3 ( .A0(n23), .A1(n29), .A2(n22), .B0(n30), .B1(in[5]), .B2(in[4]), 
        .Y(n28) );
  CLKINVX40 U22 ( .A(n28), .Y(n8) );
  CLKINVX40 U23 ( .A(in[6]), .Y(n29) );
  AOI21BX4 U24 ( .A0(n24), .A1(n9), .B0N(in[6]), .Y(n30) );
endmodule


module total_3_test_5 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n62, n63, w5_4_, n8, n9, n10, n51, n52, n53, n54, n55, n56, n57, n58,
         n61;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_171 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_170 sm_tc_2 ( .out(b1), .in({b[4:2], n61, b[0]}) );
  sm_tc_169 sm_tc_3 ( .out(c1), .in({n8, c[3:0]}) );
  sm_tc_168 sm_tc_4 ( .out(in1), .in(in) );
  add_42 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_171 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_170 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_169 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_168 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n57), .CK(clk), .RN(n9), .Q(
        up1[0]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n58), .CK(clk), .RN(n9), 
        .Q(up3[4]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n54), .CK(clk), .RN(n10), 
        .Q(h) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n53), .CK(clk), .RN(n9), 
        .Q(n63) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n55), .CK(clk), .RN(n9), 
        .Q(up3[2]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n57), .CK(clk), .RN(n10), 
        .Q(up1[3]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n53), .CK(clk), .RN(n9), 
        .Q(up3[0]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n52), .CK(clk), .RN(n9), 
        .Q(up2[0]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n55), .CK(clk), .RN(n9), 
        .Q(up2[4]) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n54), .CK(clk), .RN(n10), 
        .Q(up1[4]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n54), .CK(clk), .RN(n9), 
        .Q(up3[1]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n52), .CK(clk), .RN(n9), 
        .Q(n62) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n55), .CK(clk), .RN(n9), 
        .Q(up2[2]) );
  BUFX2 U3 ( .A(c[4]), .Y(n8) );
  CLKBUFX1TH U4 ( .A(rst), .Y(n10) );
  CLKBUFX4TH U5 ( .A(rst), .Y(n9) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n54), .CK(clk), .RN(n9), 
        .Q(up2[1]) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n55), .CK(clk), .RN(n9), 
        .Q(up1[1]) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n58), .CK(clk), .RN(n9), 
        .Q(up1[2]) );
  DLY1X1TH U38 ( .A(n56), .Y(n51) );
  INVXLTH U39 ( .A(n51), .Y(n52) );
  INVXLTH U40 ( .A(n51), .Y(n53) );
  DLY1X1TH U41 ( .A(test_se), .Y(n54) );
  DLY1X1TH U42 ( .A(test_se), .Y(n55) );
  INVXLTH U43 ( .A(test_se), .Y(n56) );
  INVXLTH U44 ( .A(n51), .Y(n57) );
  INVXLTH U45 ( .A(n51), .Y(n58) );
  DLY1X1TH U46 ( .A(n63), .Y(up3[3]) );
  DLY1X1TH U47 ( .A(n62), .Y(up2[3]) );
  CLKBUFX40 U48 ( .A(b[1]), .Y(n61) );
endmodule


module sm_tc_167 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n21, n22, n23, n28, n29, n32, n33;

  OAI2BB2X2 U2 ( .B0(n29), .B1(n6), .A0N(in[1]), .A1N(n29), .Y(out[1]) );
  CLKNAND2X4TH U3 ( .A(n22), .B(n23), .Y(n4) );
  INVX1TH U4 ( .A(in[2]), .Y(n28) );
  INVX6 U6 ( .A(in[4]), .Y(n29) );
  OAI22X1TH U7 ( .A0(n33), .A1(n28), .B0(n29), .B1(n5), .Y(out[2]) );
  DLY1X1TH U8 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX1 U9 ( .A(out[4]), .Y(out[5]) );
  CLKNAND2X2 U10 ( .A(n7), .B(in[3]), .Y(n22) );
  NAND2X4 U11 ( .A(n32), .B(n21), .Y(n23) );
  AOI31X1 U12 ( .A0(n3), .A1(n4), .A2(n5), .B0(n29), .Y(out[4]) );
  OAI2BB2X1TH U13 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  CLKBUFX2TH U17 ( .A(in[0]), .Y(out[0]) );
  AO21X4 U18 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X6 U19 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX1 U20 ( .A(in[3]), .Y(n21) );
  NOR2BXLTH U21 ( .AN(n6), .B(in[0]), .Y(n3) );
  XOR2X1 U5 ( .A(in[2]), .B(n8), .Y(n5) );
  AND2X8 U14 ( .A(n8), .B(n28), .Y(n32) );
  CLKINVX40 U15 ( .A(n32), .Y(n7) );
  CLKINVX40 U16 ( .A(n29), .Y(n33) );
endmodule


module sm_tc_166 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n6, n7, n8, n18, n19, n20, n24, n25, n28, n29;

  AOI31X4 U2 ( .A0(n3), .A1(n4), .A2(n20), .B0(n29), .Y(out[4]) );
  OR2X2 U3 ( .A(n29), .B(n20), .Y(n19) );
  INVX4 U4 ( .A(in[4]), .Y(n24) );
  NOR2BX1 U5 ( .AN(n6), .B(out[0]), .Y(n3) );
  OAI2BB2X1TH U6 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  AO21X1TH U7 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X4 U8 ( .A(in[1]), .B(out[0]), .Y(n8) );
  CLKBUFX4TH U9 ( .A(in[0]), .Y(out[0]) );
  INVX1TH U10 ( .A(in[2]), .Y(n25) );
  OAI2BB2X2 U11 ( .B0(n29), .B1(n6), .A0N(in[1]), .A1N(n29), .Y(out[1]) );
  XNOR2X2TH U12 ( .A(n7), .B(in[3]), .Y(n4) );
  OR2X2 U13 ( .A(in[4]), .B(n25), .Y(n18) );
  NAND2X8 U14 ( .A(n18), .B(n19), .Y(out[2]) );
  XOR2X1TH U15 ( .A(in[2]), .B(n8), .Y(n20) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[6]) );
  NAND2XLTH U18 ( .A(n8), .B(n25), .Y(n7) );
  CLKINVX40 U19 ( .A(n24), .Y(n28) );
  CLKINVX40 U20 ( .A(n28), .Y(n29) );
endmodule


module sm_tc_165 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n32, n36, n37, n40, n41;

  XNOR2X2 U2 ( .A(n37), .B(n8), .Y(n5) );
  NOR2X4 U4 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX2 U5 ( .A(n32), .Y(n36) );
  AOI31X2 U6 ( .A0(n3), .A1(n4), .A2(n5), .B0(n36), .Y(out[4]) );
  BUFX2TH U7 ( .A(in[4]), .Y(n32) );
  OAI2BB2X4TH U10 ( .B0(n36), .B1(n6), .A0N(in[1]), .A1N(n36), .Y(out[1]) );
  CLKBUFX1TH U11 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X1TH U13 ( .B0(n36), .B1(n4), .A0N(in[3]), .A1N(n36), .Y(out[3]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  INVX2 U17 ( .A(in[2]), .Y(n37) );
  OAI2BB1X4 U3 ( .A0N(in[0]), .A1N(in[1]), .B0(n40), .Y(n6) );
  CLKINVX40 U8 ( .A(n8), .Y(n40) );
  OAI2B2X2 U9 ( .A1N(n32), .A0(n5), .B0(n32), .B1(n37), .Y(out[2]) );
  XOR2X1 U14 ( .A(n41), .B(in[3]), .Y(n4) );
  CLKAND2X12 U18 ( .A(n8), .B(n37), .Y(n41) );
endmodule


module sm_tc_164 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n20, n21;

  OAI2BB2X2 U5 ( .B0(n21), .B1(n6), .A0N(in[1]), .A1N(n21), .Y(out[1]) );
  CLKBUFX1TH U2 ( .A(out[4]), .Y(out[6]) );
  NOR2X2TH U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI22X1TH U4 ( .A0(in[4]), .A1(n20), .B0(n21), .B1(n5), .Y(out[2]) );
  CLKBUFX1TH U6 ( .A(in[0]), .Y(out[0]) );
  AOI31X2 U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n21), .Y(out[4]) );
  NAND2XLTH U8 ( .A(n8), .B(n20), .Y(n7) );
  XNOR2X1TH U9 ( .A(n20), .B(n8), .Y(n5) );
  CLKINVX1TH U10 ( .A(in[2]), .Y(n20) );
  CLKINVX2TH U11 ( .A(in[4]), .Y(n21) );
  OAI2BB2X1TH U12 ( .B0(n21), .B1(n4), .A0N(in[3]), .A1N(n21), .Y(out[3]) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  AO21XLTH U15 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  XNOR2X1TH U16 ( .A(n7), .B(in[3]), .Y(n4) );
endmodule


module add_41_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR2X2 U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1TH U3 ( .A(B[6]), .B(A[6]), .Y(n2) );
  CLKXOR2X1TH U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_41_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n9, n1, n2, n3, n4, n5, n6, n7;
  wire   [5:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n5), .CO(carry[2]), .S(SUM[1]) );
  ADDFX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND3X4 U1 ( .A(n2), .B(n3), .C(n4), .Y(n6) );
  CLKNAND2X2 U2 ( .A(carry[5]), .B(B[5]), .Y(n3) );
  XOR2X3TH U3 ( .A(n1), .B(carry[5]), .Y(SUM[5]) );
  CLKAND2X2TH U4 ( .A(B[0]), .B(A[0]), .Y(n5) );
  CLKNAND2X2 U5 ( .A(A[5]), .B(B[5]), .Y(n4) );
  CLKXOR2X1TH U6 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X2TH U7 ( .A(B[5]), .B(A[5]), .Y(n1) );
  NAND2X1 U8 ( .A(carry[5]), .B(A[5]), .Y(n2) );
  XNOR3X4 U9 ( .A(A[6]), .B(B[6]), .C(n6), .Y(n9) );
  CLKINVX40 U10 ( .A(n9), .Y(n7) );
  CLKINVX40 U11 ( .A(n7), .Y(SUM[6]) );
endmodule


module add_41_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX4TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CLKAND2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_41_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(n2), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKINVX40 U4 ( .A(A[6]), .Y(n2) );
endmodule


module add_41_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [6:2] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKNAND2X2TH U4 ( .A(B[5]), .B(A[5]), .Y(n4) );
  CLKNAND2X2 U5 ( .A(carry[5]), .B(B[5]), .Y(n2) );
  NAND3X2TH U6 ( .A(n2), .B(n3), .C(n4), .Y(carry[6]) );
  AND2X8 U1 ( .A(carry[5]), .B(A[5]), .Y(n5) );
  CLKINVX40 U7 ( .A(n5), .Y(n3) );
  XNOR3X2 U8 ( .A(carry[5]), .B(B[5]), .C(A[5]), .Y(n6) );
  CLKINVX40 U9 ( .A(n6), .Y(SUM[5]) );
endmodule


module add_41_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_41 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n16, n17, n18, n19, n20, n21, n22;

  add_41_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n22, temp1_0_}), .B({in2[6:5], n19, in2[3], n20, in2[1:0]}), 
        .SUM(out3) );
  add_41_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, n16, temp2_0_}), .B(in), .SUM(out1) );
  add_41_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n22, temp1_0_}), .B({in3[6:3], n21, in3[1:0]}), .SUM(out2)
         );
  add_41_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n22, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_41_DW01_add_4 add_30 ( .A({in2[6:5], n18, in2[3], n20, in2[1:0]}), .B({
        in3[6:3], n21, in3[1:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_41_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX1TH U1 ( .A(temp2_1_), .Y(n16) );
  BUFX2TH U2 ( .A(in3[2]), .Y(n21) );
  INVXLTH U3 ( .A(in2[4]), .Y(n17) );
  BUFX10 U4 ( .A(in2[2]), .Y(n20) );
  INVXLTH U5 ( .A(n17), .Y(n18) );
  INVXLTH U6 ( .A(n17), .Y(n19) );
  CLKBUFX40 U13 ( .A(temp1_1_), .Y(n22) );
endmodule


module tc_sm_167 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n23, n25, n26, n27, n28, n29, n30;

  BUFX4 U3 ( .A(in[6]), .Y(n23) );
  BUFX2 U4 ( .A(n23), .Y(out[4]) );
  NOR3X1TH U5 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U6 ( .A(in[1]), .Y(n30) );
  XNOR2XLTH U7 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U8 ( .A(in[2]), .Y(n29) );
  XNOR2XLTH U9 ( .A(n29), .B(n11), .Y(n10) );
  NOR2XLTH U10 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U11 ( .A(n23), .Y(n25) );
  OAI33X4TH U12 ( .A0(in[4]), .A1(n23), .A2(in[5]), .B0(n13), .B1(n26), .B2(
        n27), .Y(n8) );
  INVXLTH U13 ( .A(in[4]), .Y(n27) );
  INVXLTH U14 ( .A(in[5]), .Y(n26) );
  CLKINVX1TH U15 ( .A(in[3]), .Y(n28) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U17 ( .A0(n25), .A1(n12), .B0(n23), .B1(n30), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U18 ( .A0(n25), .A1(n10), .B0(n23), .B1(n29), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U19 ( .A0(n9), .A1(n28), .B0(n23), .Y(n7) );
  OAI211XLTH U20 ( .A0(n23), .A1(n28), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U21 ( .A0N(n28), .A1N(n9), .B0(n23), .Y(n13) );
endmodule


module tc_sm_166 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n7, n8, n9, n10, n11, n12, n13, n35, n36, n37, n38, n39, n42, n43,
         n44, n45, n47, n48, n49, n50;

  NAND3XL U3 ( .A(n38), .B(n39), .C(n10), .Y(out[2]) );
  NOR3X1 U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  INVX5 U6 ( .A(in[6]), .Y(n42) );
  AOI31X4 U11 ( .A0(in[4]), .A1(n13), .A2(in[5]), .B0(n42), .Y(n8) );
  NOR3X6 U12 ( .A(in[5]), .B(in[6]), .C(in[4]), .Y(n5) );
  OR2XLTH U13 ( .A(in[6]), .B(n45), .Y(n37) );
  OR2XLTH U14 ( .A(n42), .B(n12), .Y(n36) );
  INVX1TH U15 ( .A(in[1]), .Y(n45) );
  OR2XLTH U17 ( .A(n42), .B(n9), .Y(n38) );
  OR2XLTH U18 ( .A(in[6]), .B(n44), .Y(n39) );
  CLKINVX1TH U19 ( .A(in[3]), .Y(n43) );
  NAND2XLTH U20 ( .A(n43), .B(n7), .Y(n13) );
  XOR2XLTH U21 ( .A(in[0]), .B(n45), .Y(n12) );
  CLKBUFX1TH U22 ( .A(in[6]), .Y(out[4]) );
  NOR2XLTH U23 ( .A(in[0]), .B(in[1]), .Y(n11) );
  NAND2BXLTH U24 ( .AN(in[0]), .B(n10), .Y(out[0]) );
  INVXLTH U25 ( .A(in[2]), .Y(n44) );
  XOR2XLTH U26 ( .A(in[2]), .B(n11), .Y(n9) );
  OR4X8 U5 ( .A(n7), .B(n42), .C(n8), .D(n43), .Y(n47) );
  AOI21BX4 U7 ( .A0(n5), .A1(n43), .B0N(n47), .Y(out[3]) );
  NAND2X8 U8 ( .A(n36), .B(n37), .Y(n48) );
  CLKINVX40 U9 ( .A(n48), .Y(n35) );
  AND2X8 U10 ( .A(n10), .B(n35), .Y(n49) );
  CLKINVX40 U16 ( .A(n49), .Y(out[1]) );
  OAI21BX4 U27 ( .A0(in[6]), .A1(n5), .B0N(n8), .Y(n50) );
  CLKINVX40 U28 ( .A(n50), .Y(n10) );
endmodule


module tc_sm_165 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n23, n24, n25, n27, n28, n29, n30,
         n31, n32;

  OAI211X1TH U6 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221XL U7 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[1])
         );
  OAI221XL U8 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[2])
         );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n23) );
  INVXLTH U12 ( .A(in[6]), .Y(n20) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  OAI21XLTH U14 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U16 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U18 ( .A(in[2]), .Y(n24) );
  INVXLTH U19 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U21 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U3 ( .A(n29), .Y(n27) );
  AOI33X4 U4 ( .A0(n29), .A1(n30), .A2(n31), .B0(n32), .B1(in[5]), .B2(n27), 
        .Y(n28) );
  CLKINVX40 U5 ( .A(n28), .Y(n8) );
  CLKINVX40 U9 ( .A(in[4]), .Y(n29) );
  CLKINVX40 U10 ( .A(in[6]), .Y(n30) );
  CLKINVX40 U22 ( .A(in[5]), .Y(n31) );
  AOI21BX4 U23 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n32) );
endmodule


module tc_sm_164 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n19, n20, n22, n23, n24, n25, n26,
         n27, n29;

  INVXLTH U3 ( .A(out[4]), .Y(n22) );
  OAI221X2 U4 ( .A0(n22), .A1(n12), .B0(out[4]), .B1(n27), .C0(n20), .Y(out[1]) );
  OAI221X2 U5 ( .A0(n22), .A1(n10), .B0(out[4]), .B1(n26), .C0(n20), .Y(out[2]) );
  OAI211X2 U6 ( .A0(out[4]), .A1(n25), .B0(n7), .C0(n20), .Y(out[3]) );
  OAI33X4 U7 ( .A0(in[4]), .A1(out[4]), .A2(n29), .B0(n13), .B1(n23), .B2(n24), 
        .Y(n8) );
  BUFX8 U8 ( .A(in[6]), .Y(out[4]) );
  INVX6 U9 ( .A(n8), .Y(n19) );
  CLKINVX16 U10 ( .A(n19), .Y(n20) );
  NAND2BX1 U11 ( .AN(in[0]), .B(n20), .Y(out[0]) );
  OAI2BB1X2 U12 ( .A0N(n25), .A1N(n9), .B0(in[6]), .Y(n13) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n25) );
  INVXLTH U14 ( .A(in[4]), .Y(n24) );
  INVXLTH U15 ( .A(n29), .Y(n23) );
  XNOR2XLTH U16 ( .A(n26), .B(n11), .Y(n10) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U18 ( .A(in[2]), .Y(n26) );
  INVXLTH U19 ( .A(in[1]), .Y(n27) );
  XNOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U21 ( .A0(n9), .A1(n25), .B0(out[4]), .Y(n7) );
  NOR3X1TH U22 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX40 U23 ( .A(in[5]), .Y(n29) );
endmodule


module total_3_test_6 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n57, n58, w5_4_, n7, n8, n9, n10, n46, n47, n48, n49, n50, n51, n52,
         n53;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_167 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_166 sm_tc_2 ( .out(b1), .in({n8, b[3:0]}) );
  sm_tc_165 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_164 sm_tc_4 ( .out(in1), .in(in) );
  add_41 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2({b1[6:2], n7, b1[0]}), .in3(c1), .in(in1) );
  tc_sm_167 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_166 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_165 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_164 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n52), .CK(clk), .RN(n10), .Q(
        up1[0]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n49), .CK(clk), .RN(n9), 
        .Q(up3[3]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n47), .CK(clk), .RN(n9), 
        .Q(up1[3]) );
  SDFFRQXLTH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n49), .CK(clk), .RN(n10), 
        .Q(up1[4]) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n49), .CK(clk), .RN(n9), 
        .Q(n58) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n50), .CK(clk), .RN(n10), 
        .Q(h) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n53), .CK(clk), .RN(n9), 
        .Q(up3[2]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n53), .CK(clk), .RN(n9), 
        .Q(up2[0]) );
  SDFFRQX1TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n49), .CK(clk), .RN(n9), 
        .Q(up3[4]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n47), .CK(clk), .RN(n9), 
        .Q(up3[1]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n50), .CK(clk), .RN(n9), 
        .Q(up3[0]) );
  SDFFRQXLTH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n50), .CK(clk), .RN(n9), 
        .Q(up2[1]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n52), .CK(clk), .RN(n9), 
        .Q(up2[2]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n48), .CK(clk), .RN(n9), 
        .Q(up2[3]) );
  SDFFRQXLTH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n48), .CK(clk), .RN(n9), 
        .Q(n57) );
  CLKBUFX2 U3 ( .A(b1[1]), .Y(n7) );
  CLKBUFX1TH U4 ( .A(b[4]), .Y(n8) );
  CLKBUFX4TH U5 ( .A(rst), .Y(n9) );
  CLKBUFX1TH U6 ( .A(rst), .Y(n10) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n50), .CK(clk), .RN(n9), 
        .Q(up1[2]) );
  DLY1X1TH U39 ( .A(n57), .Y(up1[1]) );
  DLY1X1TH U40 ( .A(n51), .Y(n46) );
  INVXLTH U41 ( .A(n46), .Y(n47) );
  INVXLTH U42 ( .A(n46), .Y(n48) );
  DLY1X1TH U43 ( .A(test_se), .Y(n49) );
  DLY1X1TH U44 ( .A(test_se), .Y(n50) );
  INVXLTH U45 ( .A(test_se), .Y(n51) );
  INVXLTH U46 ( .A(n46), .Y(n52) );
  INVXLTH U47 ( .A(n46), .Y(n53) );
  DLY1X1TH U48 ( .A(n58), .Y(up2[4]) );
endmodule


module sm_tc_163 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n23, n26;

  INVX8 U2 ( .A(in[4]), .Y(n22) );
  OAI2BB2X2 U3 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  XNOR2X2 U4 ( .A(n7), .B(in[3]), .Y(n4) );
  AO21X2 U5 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  AOI31X1 U6 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  XNOR2X2 U7 ( .A(n23), .B(n8), .Y(n5) );
  BUFX2TH U8 ( .A(in[0]), .Y(out[0]) );
  CLKINVX1TH U9 ( .A(in[2]), .Y(n23) );
  NAND2XLTH U10 ( .A(n8), .B(n23), .Y(n7) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2XLTH U13 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  NOR2X6 U16 ( .A(in[1]), .B(in[0]), .Y(n8) );
  AO2B2BX4 U14 ( .A0(n22), .A1N(n23), .B0(n26), .B1N(n5), .Y(out[2]) );
  CLKINVX40 U17 ( .A(n22), .Y(n26) );
endmodule


module sm_tc_162 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n21, n22, n25;

  NOR2X8 U2 ( .A(in[1]), .B(out[0]), .Y(n8) );
  OAI2BB2X2 U3 ( .B0(n21), .B1(n6), .A0N(in[1]), .A1N(n21), .Y(out[1]) );
  OAI22X1 U4 ( .A0(in[4]), .A1(n22), .B0(n5), .B1(n21), .Y(out[2]) );
  CLKBUFX3TH U5 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1 U6 ( .A(n22), .B(n8), .Y(n5) );
  INVX2TH U7 ( .A(in[4]), .Y(n21) );
  OAI2BB2X2 U9 ( .B0(n21), .B1(n4), .A0N(in[3]), .A1N(n21), .Y(out[3]) );
  INVX1TH U11 ( .A(in[2]), .Y(n22) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[6]) );
  AOI31X2 U13 ( .A0(n3), .A1(n4), .A2(n5), .B0(n21), .Y(out[4]) );
  AO21X1 U14 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2BXLTH U15 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  XOR2X1 U8 ( .A(n25), .B(in[3]), .Y(n4) );
  CLKAND2X12 U10 ( .A(n8), .B(n22), .Y(n25) );
endmodule


module sm_tc_161 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n28, n3, n4, n5, n6, n7, n8, n17, n19, n22, n23, n26;

  NOR2BX1 U2 ( .AN(n6), .B(in[0]), .Y(n3) );
  NOR2X2 U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX3TH U4 ( .A(in[4]), .Y(n23) );
  OAI22X2 U5 ( .A0(n17), .A1(n22), .B0(n23), .B1(n5), .Y(out[2]) );
  XNOR2X2TH U6 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2X1TH U7 ( .A(n8), .B(n22), .Y(n7) );
  INVX1TH U8 ( .A(out[4]), .Y(n19) );
  OAI2BB2X1TH U9 ( .B0(n23), .B1(n4), .A0N(in[3]), .A1N(n23), .Y(out[3]) );
  INVX1TH U10 ( .A(in[2]), .Y(n22) );
  AO21X2TH U11 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2X2TH U12 ( .B0(n23), .B1(n6), .A0N(in[1]), .A1N(n23), .Y(out[1]) );
  CLKBUFX2TH U13 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U14 ( .A(n23), .Y(n17) );
  AOI31X2TH U15 ( .A0(n3), .A1(n4), .A2(n5), .B0(n23), .Y(n28) );
  XNOR2X1TH U16 ( .A(n22), .B(n8), .Y(n5) );
  INVXLTH U17 ( .A(n19), .Y(out[5]) );
  INVXLTH U18 ( .A(n19), .Y(out[6]) );
  CLKINVX40 U19 ( .A(n28), .Y(n26) );
  CLKINVX40 U20 ( .A(n26), .Y(out[4]) );
endmodule


module sm_tc_160 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  CLKBUFX1TH U2 ( .A(in[0]), .Y(out[0]) );
  NAND2X1TH U3 ( .A(n8), .B(n21), .Y(n7) );
  XNOR2X1TH U4 ( .A(n7), .B(in[3]), .Y(n4) );
  NOR2X2TH U5 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVXLTH U6 ( .A(n18), .Y(out[6]) );
  OAI2BB2X1TH U7 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  OAI22X2TH U8 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  CLKINVX1TH U9 ( .A(in[2]), .Y(n21) );
  OAI2BB2X1TH U10 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  INVXLTH U11 ( .A(out[4]), .Y(n18) );
  INVXLTH U12 ( .A(n18), .Y(out[5]) );
  AOI31X2TH U13 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX2TH U15 ( .A(in[4]), .Y(n22) );
  XNOR2X1TH U16 ( .A(n21), .B(n8), .Y(n5) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_40_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR3X4TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_40_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKAND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_40_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X2 U1 ( .A(B[6]), .B(A[6]), .Y(n2) );
  CLKXOR2X8 U2 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  CLKAND2X2TH U3 ( .A(A[0]), .B(B[0]), .Y(n1) );
  CLKXOR2X1TH U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_40_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n3, n4, n5, n6, n7;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  NAND2XL U1 ( .A(A[6]), .B(B[6]), .Y(n5) );
  NAND2X2 U2 ( .A(n3), .B(n4), .Y(n6) );
  NAND2X6 U3 ( .A(n5), .B(n6), .Y(n7) );
  INVX2 U4 ( .A(A[6]), .Y(n3) );
  INVXLTH U5 ( .A(B[6]), .Y(n4) );
  XNOR2X4 U6 ( .A(n7), .B(carry[6]), .Y(SUM[6]) );
  AND2XLTH U7 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U8 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_40_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHX4TH U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_40_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_40 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n24, n25, n26, n27, n28;

  add_40_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n28, temp1_2_, 
        temp1_1_, n27}), .B({in2[6:3], n25, in2[1:0]}), .SUM(out3) );
  add_40_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B({in[6:2], n24, in[0]}), .SUM(out1)
         );
  add_40_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n28, temp1_2_, 
        temp1_1_, n27}), .B({in3[6:2], n26, in3[0]}), .SUM(out2) );
  add_40_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n28, temp1_2_, 
        temp1_1_, n27}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_40_DW01_add_4 add_30 ( .A({in2[6:3], n25, in2[1:0]}), .B({in3[6:2], n26, 
        in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_40_DW01_add_5 add_29 ( .A({in[6:2], n24, in[0]}), .B(in1), .SUM({
        temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_})
         );
  BUFX2 U1 ( .A(in[1]), .Y(n24) );
  CLKBUFX40 U2 ( .A(in2[2]), .Y(n25) );
  CLKBUFX40 U3 ( .A(in3[1]), .Y(n26) );
  CLKBUFX40 U4 ( .A(temp1_0_), .Y(n27) );
  CLKBUFX40 U5 ( .A(temp1_3_), .Y(n28) );
endmodule


module tc_sm_163 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n28) );
  XNOR2XLTH U7 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXLTH U10 ( .A(in[5]), .Y(n25) );
  INVXLTH U11 ( .A(in[4]), .Y(n26) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n27) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n24) );
  OAI21XLTH U16 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  OAI221XLTH U17 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U18 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(
        out[2]) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_162 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n22, n23, n24, n25, n27, n28,
         n29, n30, n31, n32;

  OAI221X1 U4 ( .A0(n29), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[1])
         );
  INVXLTH U5 ( .A(in[6]), .Y(n20) );
  OAI221X2TH U6 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[2]) );
  OAI211X1TH U7 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
  INVX2TH U8 ( .A(in[4]), .Y(n22) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U13 ( .A(n24), .B(n11), .Y(n10) );
  OAI21XLTH U14 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVX2 U16 ( .A(in[5]), .Y(n21) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U18 ( .A(in[2]), .Y(n24) );
  INVXLTH U19 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n12) );
  CLKBUFX40 U3 ( .A(n28), .Y(n27) );
  AOI33X4 U10 ( .A0(n22), .A1(n29), .A2(n21), .B0(n32), .B1(n30), .B2(n31), 
        .Y(n28) );
  CLKINVX40 U21 ( .A(n27), .Y(n8) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n29) );
  CLKINVX40 U23 ( .A(n21), .Y(n30) );
  CLKINVX40 U24 ( .A(n22), .Y(n31) );
  AOI21BX4 U25 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n32) );
endmodule


module tc_sm_161 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n18, n19, n20, n22, n23, n24, n25, n26,
         n27;

  AOI33X4 U3 ( .A0(n24), .A1(n19), .A2(n23), .B0(n20), .B1(in[5]), .B2(in[4]), 
        .Y(n18) );
  CLKINVX40 U4 ( .A(n18), .Y(n8) );
  CLKINVX40 U5 ( .A(in[6]), .Y(n19) );
  AOI21BX2 U6 ( .A0(n25), .A1(n9), .B0N(in[6]), .Y(n20) );
  OAI221XL U7 ( .A0(n22), .A1(n10), .B0(in[6]), .B1(n26), .C0(n8), .Y(out[2])
         );
  OAI221XL U8 ( .A0(n22), .A1(n12), .B0(in[6]), .B1(n27), .C0(n8), .Y(out[1])
         );
  OAI211XL U9 ( .A0(in[6]), .A1(n25), .B0(n7), .C0(n8), .Y(out[3]) );
  INVXLTH U10 ( .A(in[4]), .Y(n24) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n25) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U14 ( .A(in[1]), .Y(n27) );
  XNOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U16 ( .A(n26), .B(n11), .Y(n10) );
  INVXLTH U17 ( .A(in[2]), .Y(n26) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI21XLTH U19 ( .A0(n9), .A1(n25), .B0(in[6]), .Y(n7) );
  INVX2 U20 ( .A(in[5]), .Y(n23) );
  NAND2BXLTH U21 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U22 ( .A(in[6]), .Y(n22) );
endmodule


module tc_sm_160 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n20, n21, n22, n23, n25;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  INVX2TH U3 ( .A(in[6]), .Y(n20) );
  AOI2BB1X4 U5 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  NOR3X1TH U6 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U8 ( .A(in[6]), .Y(out[4]) );
  XOR2XLTH U9 ( .A(in[0]), .B(n23), .Y(n10) );
  INVXLTH U10 ( .A(in[1]), .Y(n23) );
  INVXLTH U11 ( .A(in[2]), .Y(n22) );
  XOR2XLTH U12 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI21XLTH U14 ( .A0(n7), .A1(n21), .B0(in[6]), .Y(n5) );
  OAI211XLTH U15 ( .A0(in[6]), .A1(n21), .B0(n5), .C0(n6), .Y(out[3]) );
  INVXLTH U16 ( .A(in[3]), .Y(n21) );
  OAI221XLTH U17 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n23), .C0(n6), .Y(
        out[1]) );
  OAI221XLTH U18 ( .A0(n20), .A1(n8), .B0(in[6]), .B1(n22), .C0(n6), .Y(out[2]) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  AO21X4 U4 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n25) );
  CLKINVX40 U20 ( .A(n25), .Y(n6) );
endmodule


module total_3_test_7 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n58, w5_4_, n5, n6, n46, n47, n48, n49, n50, n51, n52, n53;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_163 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_162 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_161 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_160 sm_tc_4 ( .out(in1), .in(in) );
  add_40 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_163 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_162 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_161 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_160 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n49), .CK(clk), .RN(n6), .Q(
        h) );
  SDFFRQXLTH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n48), .CK(clk), .RN(n5), .Q(
        up1[0]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n52), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRQX1TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n47), .CK(clk), .RN(n6), 
        .Q(up3[4]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n47), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n53), .CK(clk), .RN(n5), 
        .Q(up1[2]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(n58) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up2[1]) );
  SDFFRQX2 up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n53), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQX2 up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n52), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n6) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n5) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRX4 up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up3[3]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(up1[3]) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  DLY1X1TH U37 ( .A(n58), .Y(up2[2]) );
  DLY1X1TH U38 ( .A(n51), .Y(n46) );
  INVXLTH U39 ( .A(n46), .Y(n47) );
  INVXLTH U40 ( .A(n46), .Y(n48) );
  DLY1X1TH U41 ( .A(test_se), .Y(n49) );
  DLY1X1TH U42 ( .A(test_se), .Y(n50) );
  INVXLTH U43 ( .A(test_se), .Y(n51) );
  INVXLTH U44 ( .A(n46), .Y(n52) );
  INVXLTH U45 ( .A(n46), .Y(n53) );
endmodule


module sm_tc_159 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n21, n22;

  XNOR2X1 U2 ( .A(n7), .B(in[3]), .Y(n4) );
  BUFX2 U3 ( .A(in[4]), .Y(n17) );
  NOR2X3 U4 ( .A(in[1]), .B(out[0]), .Y(n8) );
  BUFX4 U5 ( .A(in[0]), .Y(out[0]) );
  AO21X2 U6 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NAND2XLTH U7 ( .A(n8), .B(n21), .Y(n7) );
  OAI22XLTH U8 ( .A0(n17), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  XNOR2X1 U9 ( .A(n21), .B(n8), .Y(n5) );
  INVX1TH U10 ( .A(in[2]), .Y(n21) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2XLTH U12 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  AOI31X2TH U13 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2X2TH U15 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVX4 U17 ( .A(n17), .Y(n22) );
endmodule


module sm_tc_158 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n17, n19, n22, n23, n26;

  INVX6 U2 ( .A(in[4]), .Y(n22) );
  BUFX10 U3 ( .A(in[0]), .Y(n17) );
  CLKINVX8 U4 ( .A(out[4]), .Y(n19) );
  AOI31X2 U5 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  OAI22XL U6 ( .A0(in[4]), .A1(n23), .B0(n22), .B1(n5), .Y(out[2]) );
  XNOR2X1 U7 ( .A(n23), .B(n8), .Y(n5) );
  NOR2X4 U9 ( .A(in[1]), .B(n17), .Y(n8) );
  OAI2BB2X2 U10 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  AO21X4 U11 ( .A0(n17), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKBUFX2TH U12 ( .A(n17), .Y(out[0]) );
  OAI2BB2X1TH U13 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  INVXLTH U14 ( .A(n19), .Y(out[5]) );
  INVXLTH U15 ( .A(n19), .Y(out[6]) );
  INVX2 U17 ( .A(in[2]), .Y(n23) );
  NOR2BXLTH U18 ( .AN(n6), .B(n17), .Y(n3) );
  XOR2X1 U8 ( .A(n26), .B(in[3]), .Y(n4) );
  CLKAND2X12 U16 ( .A(n8), .B(n23), .Y(n26) );
endmodule


module sm_tc_157 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n30, n31, n33, n34, n35;

  CLKBUFX3 U2 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1 U3 ( .A(n31), .B(n8), .Y(n5) );
  NOR2X2 U4 ( .A(in[1]), .B(out[0]), .Y(n8) );
  INVX1TH U5 ( .A(in[2]), .Y(n31) );
  INVX2TH U6 ( .A(in[4]), .Y(n30) );
  AOI31X2 U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n34), .Y(out[6]) );
  OAI22X1 U9 ( .A0(in[4]), .A1(n31), .B0(n34), .B1(n5), .Y(out[2]) );
  OAI2BB2X1TH U10 ( .B0(n34), .B1(n4), .A0N(in[3]), .A1N(n34), .Y(out[3]) );
  XNOR2X2TH U11 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKNAND2X2 U12 ( .A(n8), .B(n31), .Y(n7) );
  NOR2BXLTH U13 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[6]), .Y(out[4]) );
  CLKBUFX1TH U15 ( .A(out[6]), .Y(out[5]) );
  AO21X2 U16 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKINVX40 U8 ( .A(n30), .Y(n33) );
  CLKINVX40 U17 ( .A(n33), .Y(n34) );
  AO2B2X4 U18 ( .B0(in[1]), .B1(n34), .A0(n35), .A1N(n34), .Y(out[1]) );
  CLKINVX40 U19 ( .A(n6), .Y(n35) );
endmodule


module sm_tc_156 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  NOR2X2 U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI2BB2X1TH U3 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U4 ( .A(in[0]), .Y(out[0]) );
  AOI31X2TH U5 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  XNOR2X2TH U6 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI22X1TH U7 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  OAI2BB2X1TH U8 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  INVXLTH U9 ( .A(n18), .Y(out[6]) );
  CLKINVX1TH U10 ( .A(in[2]), .Y(n21) );
  CLKINVX2TH U11 ( .A(in[4]), .Y(n22) );
  INVXLTH U12 ( .A(out[4]), .Y(n18) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U14 ( .A(n18), .Y(out[5]) );
  XNOR2X1TH U15 ( .A(n21), .B(n8), .Y(n5) );
  NAND2XLTH U16 ( .A(n8), .B(n21), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_39_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX2TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX4TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X4 U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U3 ( .A(B[6]), .B(A[6]), .Y(n2) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_39_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_39_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4;
  wire   [6:2] carry;

  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR2X4 U3 ( .A(A[6]), .B(B[6]), .Y(n2) );
  XNOR2X4 U4 ( .A(carry[6]), .B(n3), .Y(n4) );
  CLKINVX20 U5 ( .A(n2), .Y(n3) );
  CLKINVX40 U6 ( .A(n4), .Y(SUM[6]) );
endmodule


module add_39_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_39_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n3, n4, n5, n6, n7;
  wire   [6:2] carry;

  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n5), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  NAND2X2TH U1 ( .A(n3), .B(n4), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n5) );
  NAND2XLTH U3 ( .A(B[0]), .B(n7), .Y(n3) );
  INVXLTH U4 ( .A(B[0]), .Y(n6) );
  INVXLTH U5 ( .A(A[0]), .Y(n7) );
  NAND2XLTH U6 ( .A(n6), .B(A[0]), .Y(n4) );
endmodule


module add_39_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n3, n1;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2TH U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(n3) );
  ADDFX2TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(carry[3]), .CI(B[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKBUFX40 U3 ( .A(n3), .Y(SUM[2]) );
endmodule


module add_39 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n18, n19, n20, n21, n22, n23, n24;

  add_39_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n23, n18}), .B({in2[6:1], n22}), .SUM(out3) );
  add_39_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, n20}), .B({in[6:2], n19, in[0]}), .SUM(out1) );
  add_39_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, n18}), .B({n21, in3[5:1], n24}), .SUM(out2) );
  add_39_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n23, n18}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_39_DW01_add_4 add_30 ( .A({in2[6:1], n22}), .B({n21, in3[5:1], n24}), 
        .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, 
        temp2_0_}) );
  add_39_DW01_add_5 add_29 ( .A({in[6:2], n19, in[0]}), .B(in1), .SUM({
        temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_})
         );
  BUFX2TH U1 ( .A(in[1]), .Y(n19) );
  BUFX2 U2 ( .A(temp1_0_), .Y(n18) );
  BUFX3TH U3 ( .A(temp2_0_), .Y(n20) );
  CLKBUFX1TH U4 ( .A(in3[6]), .Y(n21) );
  CLKBUFX40 U5 ( .A(in2[0]), .Y(n22) );
  CLKBUFX40 U6 ( .A(temp1_1_), .Y(n23) );
  CLKBUFX40 U13 ( .A(in3[0]), .Y(n24) );
endmodule


module tc_sm_159 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n25, n26, n28, n29, n30, n31, n32;

  CLKINVX1TH U3 ( .A(n25), .Y(n26) );
  CLKINVX1TH U4 ( .A(in[6]), .Y(n25) );
  CLKBUFX1TH U5 ( .A(in[6]), .Y(out[4]) );
  NOR3X1TH U6 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U7 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U9 ( .A(in[2]), .Y(n31) );
  XNOR2XLTH U10 ( .A(n31), .B(n11), .Y(n10) );
  NOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U12 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n28), .B2(
        n29), .Y(n8) );
  INVXLTH U13 ( .A(in[5]), .Y(n28) );
  INVXLTH U14 ( .A(in[4]), .Y(n29) );
  CLKINVX1TH U15 ( .A(in[3]), .Y(n30) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U17 ( .A0(n25), .A1(n12), .B0(n26), .B1(n32), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U18 ( .A0(n25), .A1(n10), .B0(n26), .B1(n31), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U19 ( .A0(n9), .A1(n30), .B0(in[6]), .Y(n7) );
  OAI211XLTH U20 ( .A0(n26), .A1(n30), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U21 ( .A0N(n30), .A1N(n9), .B0(n26), .Y(n13) );
endmodule


module tc_sm_158 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n25, n27, n28, n29, n30;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OAI221X1 U3 ( .A0(n27), .A1(n8), .B0(in[6]), .B1(n29), .C0(n6), .Y(out[2])
         );
  OAI211XL U4 ( .A0(in[6]), .A1(n28), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI221XL U5 ( .A0(n27), .A1(n10), .B0(in[6]), .B1(n30), .C0(n6), .Y(out[1])
         );
  OAI21BX2TH U6 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n25) );
  AOI21BX4 U8 ( .A0(in[6]), .A1(n11), .B0N(n25), .Y(n6) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  XOR2XLTH U10 ( .A(in[0]), .B(n30), .Y(n10) );
  INVXLTH U11 ( .A(in[1]), .Y(n30) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI21XLTH U13 ( .A0(n7), .A1(n28), .B0(in[6]), .Y(n5) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U15 ( .A(in[6]), .Y(n27) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  INVXLTH U17 ( .A(in[3]), .Y(n28) );
  INVXLTH U18 ( .A(in[2]), .Y(n29) );
  XOR2XLTH U19 ( .A(in[2]), .B(n9), .Y(n8) );
endmodule


module tc_sm_157 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n18, n19, n20, n22, n23, n24, n25, n26,
         n27;

  CLKINVX12 U3 ( .A(n18), .Y(n8) );
  INVXLTH U4 ( .A(in[5]), .Y(n23) );
  INVXLTH U5 ( .A(in[6]), .Y(n22) );
  NOR3X1TH U6 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U7 ( .A(in[3]), .Y(n25) );
  INVXLTH U8 ( .A(in[4]), .Y(n24) );
  AOI21BXLTH U9 ( .A0(n25), .A1(n9), .B0N(in[6]), .Y(n20) );
  INVXLTH U10 ( .A(in[6]), .Y(n19) );
  CLKBUFX1TH U11 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U12 ( .A(n26), .B(n11), .Y(n10) );
  NOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI21XLTH U14 ( .A0(n9), .A1(n25), .B0(in[6]), .Y(n7) );
  INVXLTH U15 ( .A(in[1]), .Y(n27) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  AOI33X4 U17 ( .A0(n24), .A1(n19), .A2(n23), .B0(n20), .B1(in[5]), .B2(in[4]), 
        .Y(n18) );
  OAI221XLTH U18 ( .A0(n22), .A1(n12), .B0(in[6]), .B1(n27), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U19 ( .A0(n22), .A1(n10), .B0(in[6]), .B1(n26), .C0(n8), .Y(
        out[2]) );
  INVXLTH U20 ( .A(in[2]), .Y(n26) );
  NAND2BXLTH U21 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211XLTH U22 ( .A0(in[6]), .A1(n25), .B0(n7), .C0(n8), .Y(out[3]) );
endmodule


module tc_sm_156 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n19, n20, n21, n22, n23, n24, n26,
         n27;

  OAI2BB1X4 U3 ( .A0N(n22), .A1N(n9), .B0(in[6]), .Y(n13) );
  NAND2BX1TH U4 ( .AN(in[0]), .B(n27), .Y(out[0]) );
  OAI211X2TH U5 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n27), .Y(out[3]) );
  INVXLTH U6 ( .A(in[6]), .Y(n19) );
  OAI221X2TH U7 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n27), .Y(
        out[1]) );
  OAI221X2TH U8 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n27), .Y(
        out[2]) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n22) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVX2TH U11 ( .A(in[4]), .Y(n21) );
  INVX2TH U12 ( .A(in[5]), .Y(n20) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U14 ( .A(n23), .B(n11), .Y(n10) );
  INVXLTH U15 ( .A(in[2]), .Y(n23) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U17 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U19 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  OAI33X4 U20 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n20), .B2(
        n21), .Y(n8) );
  CLKINVX40 U21 ( .A(n8), .Y(n26) );
  CLKINVX40 U22 ( .A(n26), .Y(n27) );
endmodule


module total_3_test_8 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n63, w5_4_, n4, n5, n6, n41, n42, n43, n52, n53, n54, n55, n56, n57,
         n58, n59;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_159 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_158 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_157 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_156 sm_tc_4 ( .out(in1), .in(in) );
  add_39 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1({a1[6:1], 
        n4}), .in2(b1), .in3(c1), .in(in1) );
  tc_sm_159 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_158 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_157 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_156 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n53), .CK(clk), .RN(n5), .Q(
        up1[0]) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n58), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n56), .CK(clk), .RN(n6), .Q(
        h) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n54), .CK(clk), .RN(n5), 
        .Q(n63) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n55), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRQX2TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n55), .CK(clk), .RN(n6), 
        .Q(up3[4]) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n59), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQX1TH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n54), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n59), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n55), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n58), .CK(clk), .RN(n6), 
        .Q(up1[2]) );
  CLKBUFX1TH U3 ( .A(a1[0]), .Y(n4) );
  CLKBUFX1TH U4 ( .A(rst), .Y(n6) );
  CLKBUFX4TH U5 ( .A(rst), .Y(n5) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n56), .CK(clk), .RN(n5), 
        .Q(up2[1]) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n56), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  SDFFRX4 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n53), .CK(clk), .RN(n5), 
        .Q(up2[2]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n55), .CK(clk), .RN(n5), 
        .Q(up1[3]) );
  SDFFRX4 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n56), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  INVXLTH U38 ( .A(test_se), .Y(n41) );
  INVXLTH U39 ( .A(n41), .Y(n42) );
  INVXLTH U40 ( .A(n41), .Y(n43) );
  DLY1X1TH U41 ( .A(n57), .Y(n52) );
  INVXLTH U42 ( .A(n52), .Y(n53) );
  INVXLTH U43 ( .A(n52), .Y(n54) );
  DLY1X1TH U44 ( .A(n42), .Y(n55) );
  DLY1X1TH U45 ( .A(n43), .Y(n56) );
  INVXLTH U46 ( .A(n42), .Y(n57) );
  INVXLTH U47 ( .A(n52), .Y(n58) );
  INVXLTH U48 ( .A(n52), .Y(n59) );
  DLY1X1TH U49 ( .A(n63), .Y(up3[3]) );
endmodule


module sm_tc_155 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n23, n26, n27, n28;

  INVX6 U3 ( .A(in[4]), .Y(n22) );
  OAI2BB2X4TH U5 ( .B0(n27), .B1(n6), .A0N(in[1]), .A1N(n27), .Y(out[1]) );
  AO21X2 U6 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X4 U7 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U8 ( .A(in[2]), .Y(n23) );
  XNOR2X4TH U9 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX1TH U10 ( .A(out[4]), .Y(out[6]) );
  OAI22X2 U11 ( .A0(in[4]), .A1(n23), .B0(n27), .B1(n5), .Y(out[2]) );
  AOI31X2TH U12 ( .A0(n3), .A1(n4), .A2(n5), .B0(n27), .Y(out[4]) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2XLTH U14 ( .B0(n27), .B1(n4), .A0N(in[3]), .A1N(n27), .Y(out[3]) );
  BUFX2TH U15 ( .A(in[0]), .Y(out[0]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX40 U2 ( .A(n22), .Y(n26) );
  CLKINVX40 U4 ( .A(n26), .Y(n27) );
  XOR2X1 U17 ( .A(in[2]), .B(n8), .Y(n5) );
  AND2X8 U18 ( .A(n8), .B(n23), .Y(n28) );
  CLKINVX40 U19 ( .A(n28), .Y(n7) );
endmodule


module sm_tc_154 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n23, n24, n25, n26, n27, n28, n29, n33;

  OAI2BB2X2 U2 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  BUFX10 U3 ( .A(in[0]), .Y(out[0]) );
  NOR2XLTH U4 ( .A(in[4]), .B(n33), .Y(n23) );
  OR2X2 U6 ( .A(n23), .B(n24), .Y(out[2]) );
  INVX6 U7 ( .A(in[4]), .Y(n29) );
  NAND2X2TH U8 ( .A(n8), .B(n33), .Y(n7) );
  NAND2X2 U9 ( .A(n27), .B(n28), .Y(n4) );
  NOR2X2 U10 ( .A(in[1]), .B(out[0]), .Y(n8) );
  CLKNAND2X2TH U11 ( .A(n25), .B(n26), .Y(n28) );
  XNOR2X1 U12 ( .A(n33), .B(n8), .Y(n5) );
  INVXLTH U13 ( .A(n7), .Y(n25) );
  AOI31X4TH U14 ( .A0(n3), .A1(n5), .A2(n4), .B0(n29), .Y(out[4]) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[6]) );
  NAND2XLTH U16 ( .A(n7), .B(in[3]), .Y(n27) );
  INVXLTH U17 ( .A(in[3]), .Y(n26) );
  AO21X2 U18 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2X1TH U19 ( .B0(n29), .B1(n6), .A0N(in[1]), .A1N(n29), .Y(out[1]) );
  CLKINVX1TH U20 ( .A(in[2]), .Y(n33) );
  NOR2BXLTH U21 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKBUFX1TH U22 ( .A(out[4]), .Y(out[5]) );
  NOR2BX8 U5 ( .AN(in[4]), .B(n5), .Y(n24) );
endmodule


module sm_tc_153 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n19, n20, n21, n25, n26;

  OAI2BB2X2 U2 ( .B0(n25), .B1(n6), .A0N(in[1]), .A1N(n25), .Y(out[1]) );
  NOR2X2 U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX4 U4 ( .A(in[4]), .Y(n25) );
  INVX2 U5 ( .A(in[2]), .Y(n26) );
  XNOR2X2 U6 ( .A(n26), .B(n8), .Y(n5) );
  AO21X2TH U7 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NAND3XL U8 ( .A(n3), .B(n4), .C(n5), .Y(n19) );
  CLKBUFX2TH U9 ( .A(out[5]), .Y(out[4]) );
  OR2XLTH U10 ( .A(n25), .B(n5), .Y(n21) );
  CLKBUFX1TH U11 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X1TH U12 ( .B0(n25), .B1(n4), .A0N(in[3]), .A1N(n25), .Y(out[3]) );
  AND2X1TH U13 ( .A(n19), .B(in[4]), .Y(out[5]) );
  CLKBUFX1TH U14 ( .A(out[5]), .Y(out[6]) );
  OR2XLTH U15 ( .A(in[4]), .B(n26), .Y(n20) );
  NAND2X1TH U16 ( .A(n20), .B(n21), .Y(out[2]) );
  XNOR2X4 U17 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U18 ( .A(n8), .B(n26), .Y(n7) );
  NOR2BXLTH U19 ( .AN(n6), .B(in[0]), .Y(n3) );
endmodule


module sm_tc_152 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n28, n31, n32;

  NOR2X4 U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  AOI31X2TH U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n32), .Y(out[4]) );
  NAND2X2 U4 ( .A(n8), .B(n31), .Y(n7) );
  INVX2 U5 ( .A(in[2]), .Y(n31) );
  NAND2X2TH U6 ( .A(n25), .B(n26), .Y(n4) );
  NAND2X2TH U7 ( .A(n23), .B(n24), .Y(n26) );
  OAI2BB2X2TH U8 ( .B0(n32), .B1(n4), .A0N(in[3]), .A1N(n32), .Y(out[3]) );
  NAND2X1TH U9 ( .A(n17), .B(n18), .Y(out[2]) );
  OR2X1TH U10 ( .A(n32), .B(n5), .Y(n18) );
  OR2XLTH U11 ( .A(in[4]), .B(n31), .Y(n17) );
  NAND2X1TH U12 ( .A(n21), .B(n22), .Y(n5) );
  NAND2XLTH U13 ( .A(n7), .B(in[3]), .Y(n25) );
  NAND2XLTH U14 ( .A(n31), .B(n8), .Y(n21) );
  NAND2XLTH U15 ( .A(n19), .B(n20), .Y(n22) );
  INVXLTH U16 ( .A(n8), .Y(n20) );
  OAI2BB2X1TH U17 ( .B0(n32), .B1(n6), .A0N(in[1]), .A1N(n32), .Y(out[1]) );
  CLKBUFX1TH U18 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U19 ( .A(n7), .Y(n23) );
  INVXLTH U20 ( .A(n31), .Y(n19) );
  INVXLTH U21 ( .A(in[3]), .Y(n24) );
  CLKINVX2TH U22 ( .A(in[4]), .Y(n32) );
  INVXLTH U23 ( .A(out[4]), .Y(n28) );
  INVXLTH U24 ( .A(n28), .Y(out[5]) );
  NOR2BXLTH U25 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U26 ( .A(n28), .Y(out[6]) );
  AO21XLTH U27 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_38_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X4TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_38_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR3X4TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_38_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_38_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n2, n3;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XNOR2X4 U1 ( .A(n3), .B(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR2XLTH U3 ( .A(A[6]), .B(B[6]), .Y(n3) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n2) );
endmodule


module add_38_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2TH U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_38_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_38 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n18, n19, n20, n21, n22;

  add_38_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in2[6:5], n20, in2[3:2], n18, 
        in2[0]}), .SUM(out3) );
  add_38_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, n22, temp2_2_, 
        temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_38_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in3[6:2], n19, n21}), .SUM(out2)
         );
  add_38_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, n22, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_38_DW01_add_4 add_30 ( .A({in2[6:5], n20, in2[3:2], n18, in2[0]}), .B({
        in3[6:2], n19, n21}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}) );
  add_38_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX6 U1 ( .A(in2[1]), .Y(n18) );
  CLKBUFX1TH U2 ( .A(in3[1]), .Y(n19) );
  CLKBUFX1TH U3 ( .A(in2[4]), .Y(n20) );
  CLKBUFX40 U4 ( .A(in3[0]), .Y(n21) );
  CLKBUFX40 U5 ( .A(temp2_3_), .Y(n22) );
endmodule


module tc_sm_155 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n28) );
  XNOR2XLTH U7 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXLTH U10 ( .A(in[4]), .Y(n26) );
  INVXLTH U11 ( .A(in[5]), .Y(n25) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n27) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n24) );
  OAI21XLTH U16 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  OAI221XLTH U17 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U18 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(
        out[2]) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_154 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n20, n21, n22, n24, n25, n26, n27,
         n28, n29;

  BUFX10 U3 ( .A(n8), .Y(n21) );
  INVX3 U4 ( .A(n22), .Y(out[4]) );
  OR2X2 U5 ( .A(n9), .B(n27), .Y(n20) );
  NAND2X2 U6 ( .A(n20), .B(out[4]), .Y(n7) );
  OAI211X1 U7 ( .A0(out[4]), .A1(n27), .B0(n7), .C0(n21), .Y(out[3]) );
  OAI221X1 U8 ( .A0(n24), .A1(n12), .B0(out[4]), .B1(n29), .C0(n21), .Y(out[1]) );
  OAI33X4 U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(n26), .Y(n8) );
  OAI2BB1X2 U10 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
  NAND2BXLTH U11 ( .AN(in[0]), .B(n21), .Y(out[0]) );
  XNOR2XLTH U12 ( .A(n28), .B(n11), .Y(n10) );
  OAI221X2TH U13 ( .A0(n24), .A1(n10), .B0(out[4]), .B1(n28), .C0(n21), .Y(
        out[2]) );
  CLKINVX1TH U14 ( .A(in[3]), .Y(n27) );
  NOR3X1TH U15 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U16 ( .A(in[4]), .Y(n26) );
  INVXLTH U17 ( .A(in[5]), .Y(n25) );
  INVXLTH U18 ( .A(in[6]), .Y(n24) );
  NOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U20 ( .A(in[2]), .Y(n28) );
  INVXLTH U21 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U22 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U23 ( .A(in[6]), .Y(n22) );
endmodule


module tc_sm_153 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n18, n19, n20, n22, n23, n24, n25, n26;

  CLKINVX4 U3 ( .A(n18), .Y(n8) );
  AOI33X4 U4 ( .A0(n23), .A1(n19), .A2(n22), .B0(n20), .B1(in[5]), .B2(in[4]), 
        .Y(n18) );
  INVX1 U5 ( .A(in[6]), .Y(n19) );
  AOI21BX2TH U6 ( .A0(n24), .A1(n9), .B0N(in[6]), .Y(n20) );
  CLKINVX1TH U7 ( .A(in[3]), .Y(n24) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U9 ( .A(in[4]), .Y(n23) );
  INVXLTH U10 ( .A(in[5]), .Y(n22) );
  NAND2BXLTH U11 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U12 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n25), .C0(n8), .Y(
        out[2]) );
  XNOR2XLTH U13 ( .A(n25), .B(n11), .Y(n10) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U15 ( .A(in[2]), .Y(n25) );
  CLKBUFX1TH U16 ( .A(in[6]), .Y(out[4]) );
  OAI221XLTH U17 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n26), .C0(n8), .Y(
        out[1]) );
  INVXLTH U18 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI211XLTH U20 ( .A0(in[6]), .A1(n24), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI21XLTH U21 ( .A0(n9), .A1(n24), .B0(in[6]), .Y(n7) );
endmodule


module tc_sm_152 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n21, n23, n24, n25, n26, n28;

  OAI211XL U3 ( .A0(in[6]), .A1(n24), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI21XL U5 ( .A0(n7), .A1(n24), .B0(in[6]), .Y(n5) );
  INVX2TH U6 ( .A(in[6]), .Y(n23) );
  AOI21BX4 U7 ( .A0(in[6]), .A1(n11), .B0N(n21), .Y(n6) );
  OAI221X2 U8 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n26), .C0(n6), .Y(out[1])
         );
  OAI221X2 U9 ( .A0(n23), .A1(n8), .B0(in[6]), .B1(n25), .C0(n6), .Y(out[2])
         );
  OAI2B11XLTH U10 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U13 ( .A(in[2]), .Y(n25) );
  XOR2XLTH U14 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n9) );
  XOR2XLTH U16 ( .A(in[0]), .B(n26), .Y(n10) );
  INVXLTH U17 ( .A(in[1]), .Y(n26) );
  INVXLTH U18 ( .A(in[3]), .Y(n24) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  AOI2BB1X4 U4 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n28) );
  CLKINVX40 U20 ( .A(n28), .Y(n21) );
endmodule


module total_3_test_9 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n56, w5_4_, n4, n5, n40, n45, n46, n47, n48, n49, n50, n51, n52;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_155 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_154 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_153 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_152 sm_tc_4 ( .out(in1), .in(in) );
  add_38 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_155 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_154 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_153 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_152 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up2[3]) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n46), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n48), .CK(clk), .RN(n5), .Q(
        h) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(n56) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRQX2TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQX1TH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up1[4]) );
  SDFFRHQX2TH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up1[1]) );
  SDFFRQX1TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up2[4]) );
  CLKBUFX4TH U3 ( .A(rst), .Y(n4) );
  CLKBUFX1TH U4 ( .A(rst), .Y(n5) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up1[2]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up1[3]) );
  SDFFRX4 up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n49), .CK(clk), .RN(n4), .Q(
        up1[0]) );
  INVXLTH U37 ( .A(n50), .Y(n40) );
  DLY1X1TH U38 ( .A(n50), .Y(n45) );
  INVXLTH U39 ( .A(n45), .Y(n46) );
  INVXLTH U40 ( .A(n45), .Y(n47) );
  DLY1X1TH U41 ( .A(n40), .Y(n48) );
  DLY1X1TH U42 ( .A(test_se), .Y(n49) );
  INVXLTH U43 ( .A(test_se), .Y(n50) );
  INVXLTH U44 ( .A(n45), .Y(n51) );
  INVXLTH U45 ( .A(n45), .Y(n52) );
  DLY1X1TH U46 ( .A(n56), .Y(up3[3]) );
endmodule


module sm_tc_151 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n21, n23, n26, n27, n30, n31;

  OAI2BB2X1 U2 ( .B0(n26), .B1(n6), .A0N(n21), .A1N(n26), .Y(out[1]) );
  INVX2 U3 ( .A(in[4]), .Y(n26) );
  INVX2TH U4 ( .A(in[2]), .Y(n27) );
  INVXLTH U5 ( .A(n23), .Y(out[6]) );
  NOR2BXLTH U6 ( .AN(n6), .B(in[0]), .Y(n3) );
  XNOR2X2TH U7 ( .A(n27), .B(n8), .Y(n5) );
  CLKBUFX1TH U8 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2XLTH U9 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  CLKBUFX1TH U10 ( .A(in[1]), .Y(n21) );
  OAI22XLTH U11 ( .A0(in[4]), .A1(n27), .B0(n26), .B1(n5), .Y(out[2]) );
  AOI31X2TH U12 ( .A0(n3), .A1(n4), .A2(n31), .B0(n26), .Y(out[4]) );
  AO21X2 U13 ( .A0(in[0]), .A1(n21), .B0(n8), .Y(n6) );
  NOR2X4 U14 ( .A(n21), .B(in[0]), .Y(n8) );
  INVXLTH U17 ( .A(out[4]), .Y(n23) );
  INVXLTH U18 ( .A(n23), .Y(out[5]) );
  XNOR2X1 U15 ( .A(n30), .B(in[3]), .Y(n4) );
  CLKNAND2X12 U16 ( .A(n8), .B(n27), .Y(n30) );
  XNOR2X2TH U19 ( .A(n27), .B(n8), .Y(n31) );
endmodule


module sm_tc_150 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n25, n26, n28, n29, n33, n34, n37;

  BUFX2 U2 ( .A(out[4]), .Y(out[5]) );
  BUFX10 U3 ( .A(in[1]), .Y(n25) );
  INVX6 U4 ( .A(in[4]), .Y(n33) );
  OAI22X1 U5 ( .A0(in[4]), .A1(n34), .B0(n33), .B1(n5), .Y(out[2]) );
  NAND2X2 U6 ( .A(n28), .B(n29), .Y(n5) );
  BUFX2TH U7 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X1 U9 ( .B0(n33), .B1(n6), .A0N(n25), .A1N(n33), .Y(out[1]) );
  INVX2TH U10 ( .A(in[2]), .Y(n34) );
  OAI2BB2XL U11 ( .B0(n33), .B1(n4), .A0N(in[3]), .A1N(n33), .Y(out[3]) );
  XNOR2X2TH U12 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U13 ( .A(n8), .B(n34), .Y(n7) );
  NAND2XLTH U14 ( .A(n26), .B(n37), .Y(n29) );
  NAND2XLTH U15 ( .A(n34), .B(n8), .Y(n28) );
  AOI31X2TH U16 ( .A0(n3), .A1(n4), .A2(n5), .B0(n33), .Y(out[4]) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  AO21X2 U18 ( .A0(in[0]), .A1(n25), .B0(n8), .Y(n6) );
  INVXL U19 ( .A(n34), .Y(n26) );
  CLKBUFX1TH U21 ( .A(out[4]), .Y(out[6]) );
  OR2X8 U8 ( .A(n25), .B(in[0]), .Y(n37) );
  CLKINVX40 U20 ( .A(n37), .Y(n8) );
endmodule


module sm_tc_149 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n23, n24, n25, n26, n30, n31;

  BUFX2TH U2 ( .A(in[0]), .Y(out[0]) );
  AO21XL U3 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X6 U4 ( .A(in[1]), .B(in[0]), .Y(n8) );
  BUFX2TH U5 ( .A(in[4]), .Y(n23) );
  INVX4 U6 ( .A(n23), .Y(n31) );
  OAI2BB2XL U7 ( .B0(n31), .B1(n4), .A0N(in[3]), .A1N(n31), .Y(out[3]) );
  XNOR2X1 U8 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI22X1 U9 ( .A0(n23), .A1(n30), .B0(n31), .B1(n5), .Y(out[2]) );
  NAND2X2 U10 ( .A(n25), .B(n26), .Y(n5) );
  INVX2TH U11 ( .A(in[2]), .Y(n30) );
  AOI31X2 U12 ( .A0(n3), .A1(n4), .A2(n5), .B0(n31), .Y(out[4]) );
  NAND2XLTH U13 ( .A(in[2]), .B(n24), .Y(n26) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X4 U16 ( .B0(n31), .B1(n6), .A0N(in[1]), .A1N(n31), .Y(out[1]) );
  NAND2XLTH U17 ( .A(n30), .B(n8), .Y(n25) );
  INVXLTH U18 ( .A(n8), .Y(n24) );
  NOR2BXLTH U19 ( .AN(n6), .B(in[0]), .Y(n3) );
  NAND2XLTH U20 ( .A(n8), .B(n30), .Y(n7) );
endmodule


module sm_tc_148 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  XNOR2X1 U2 ( .A(n21), .B(n8), .Y(n5) );
  NOR2X2TH U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X2TH U4 ( .A(n7), .B(in[3]), .Y(n4) );
  AOI31X2TH U5 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  INVXLTH U6 ( .A(out[4]), .Y(n18) );
  OAI2BB2X1TH U7 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKINVX1TH U8 ( .A(in[2]), .Y(n21) );
  NAND2XLTH U9 ( .A(n8), .B(n21), .Y(n7) );
  OAI22X1TH U10 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  CLKINVX2TH U11 ( .A(in[4]), .Y(n22) );
  NOR2BXLTH U12 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U13 ( .A(n18), .Y(out[5]) );
  INVXLTH U14 ( .A(n18), .Y(out[6]) );
  CLKBUFX1TH U15 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X2TH U16 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_37_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_37_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [6:2] carry;

  NAND2X2 U7 ( .A(n6), .B(n11), .Y(n4) );
  NAND2X2 U8 ( .A(n10), .B(carry[3]), .Y(n5) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  NAND3X2 U1 ( .A(n7), .B(n8), .C(n9), .Y(carry[4]) );
  NAND2XLTH U2 ( .A(carry[3]), .B(B[3]), .Y(n8) );
  AND2X1TH U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  INVXLTH U5 ( .A(n6), .Y(n10) );
  XOR2X1TH U6 ( .A(B[3]), .B(A[3]), .Y(n6) );
  INVXLTH U9 ( .A(carry[3]), .Y(n11) );
  NAND2XLTH U10 ( .A(A[3]), .B(B[3]), .Y(n9) );
  NAND2XLTH U11 ( .A(carry[3]), .B(A[3]), .Y(n7) );
  CLKNAND2X2 U12 ( .A(n4), .B(n5), .Y(SUM[3]) );
endmodule


module add_37_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_37_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_37_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n4, n5, n6, n7, n8, n9, n10;
  wire   [6:2] carry;

  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_2 ( .A(carry[2]), .B(A[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X2 U1 ( .A(carry[5]), .B(A[5]), .C(B[5]), .Y(SUM[5]) );
  NAND2X2 U2 ( .A(carry[5]), .B(A[5]), .Y(n6) );
  NAND2X2 U3 ( .A(carry[5]), .B(B[5]), .Y(n7) );
  NAND2XL U4 ( .A(A[5]), .B(B[5]), .Y(n8) );
  NAND3X4 U5 ( .A(n6), .B(n7), .C(n8), .Y(carry[6]) );
  NAND2X4 U6 ( .A(n4), .B(n5), .Y(SUM[0]) );
  NAND2XLTH U7 ( .A(n9), .B(A[0]), .Y(n5) );
  CLKNAND2X2TH U8 ( .A(B[0]), .B(n10), .Y(n4) );
  INVXLTH U9 ( .A(B[0]), .Y(n9) );
  INVXLTH U10 ( .A(A[0]), .Y(n10) );
  AND2XLTH U11 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_37_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2TH U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X3TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X2 U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_37 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23;

  add_37_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n23, 
        temp1_1_, temp1_0_}), .B({in2[6:5], n21, in2[3], n13, n17, n15}), 
        .SUM(out3) );
  add_37_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, n14}), .B({in[6:2], n18, in[0]}), .SUM(out1) );
  add_37_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in3[6:4], n22, in3[2:0]}), .SUM(
        out2) );
  add_37_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n23, 
        temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, n16, n19, 
        temp2_1_, n14}), .SUM(out) );
  add_37_DW01_add_4 add_30 ( .A({in2[6:3], n13, in2[1], n15}), .B({in3[6:4], 
        n22, in3[2:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}) );
  add_37_DW01_add_5 add_29 ( .A({in[6:2], n18, in[0]}), .B(in1), .SUM({
        temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_})
         );
  BUFX2 U1 ( .A(in[1]), .Y(n18) );
  DLY1X1TH U2 ( .A(in2[1]), .Y(n17) );
  BUFX6 U3 ( .A(in2[2]), .Y(n13) );
  BUFX14 U4 ( .A(temp2_0_), .Y(n14) );
  BUFX10 U5 ( .A(in2[0]), .Y(n15) );
  CLKBUFX1TH U6 ( .A(temp2_3_), .Y(n16) );
  CLKBUFX1TH U13 ( .A(temp2_2_), .Y(n19) );
  INVXLTH U14 ( .A(n20), .Y(n21) );
  INVXLTH U15 ( .A(in2[4]), .Y(n20) );
  CLKBUFX40 U16 ( .A(in3[3]), .Y(n22) );
  CLKBUFX40 U17 ( .A(temp1_2_), .Y(n23) );
endmodule


module tc_sm_151 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U10 ( .A(in[4]), .Y(n28) );
  INVXLTH U11 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_150 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n21, n22, n23, n24, n26, n27, n28,
         n29, n30, n31, n33;

  INVXLTH U3 ( .A(out[4]), .Y(n26) );
  BUFX4 U4 ( .A(n8), .Y(n22) );
  BUFX6 U5 ( .A(in[6]), .Y(out[4]) );
  NAND2X1 U7 ( .A(n22), .B(n21), .Y(out[2]) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n29) );
  OAI2BB1X4 U9 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
  INVX2 U10 ( .A(in[5]), .Y(n27) );
  OAI221XL U11 ( .A0(n26), .A1(n12), .B0(out[4]), .B1(n31), .C0(n22), .Y(
        out[1]) );
  OAI211X1TH U12 ( .A0(out[4]), .A1(n29), .B0(n7), .C0(n22), .Y(out[3]) );
  OAI33X4 U13 ( .A0(in[4]), .A1(out[4]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U14 ( .A(in[2]), .Y(n30) );
  INVX2TH U15 ( .A(in[4]), .Y(n28) );
  NOR3X1TH U16 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  OAI21XLTH U17 ( .A0(n9), .A1(n29), .B0(out[4]), .Y(n7) );
  OR2XLTH U18 ( .A(n26), .B(n10), .Y(n23) );
  XNOR2XLTH U19 ( .A(n30), .B(n11), .Y(n10) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n22), .Y(out[0]) );
  INVXLTH U21 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U22 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U23 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OR2XLTH U24 ( .A(out[4]), .B(n30), .Y(n24) );
  NAND2X8 U6 ( .A(n23), .B(n24), .Y(n33) );
  CLKINVX40 U25 ( .A(n33), .Y(n21) );
endmodule


module tc_sm_149 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n22, n23, n25, n26, n27, n29, n30, n31,
         n32, n33, n34;

  OAI211XL U3 ( .A0(n29), .A1(n25), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221XL U4 ( .A0(n22), .A1(n12), .B0(n29), .B1(n27), .C0(n8), .Y(out[1]) );
  OAI221XL U5 ( .A0(n22), .A1(n10), .B0(n29), .B1(n26), .C0(n8), .Y(out[2]) );
  INVXLTH U8 ( .A(in[6]), .Y(n22) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n25) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U12 ( .A(in[5]), .Y(n23) );
  CLKBUFX1TH U13 ( .A(n29), .Y(out[4]) );
  XNOR2XLTH U14 ( .A(n26), .B(n11), .Y(n10) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[2]), .Y(n26) );
  INVXLTH U17 ( .A(in[1]), .Y(n27) );
  XNOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U19 ( .A0(n9), .A1(n25), .B0(in[6]), .Y(n7) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  CLKINVX40 U6 ( .A(n33), .Y(n29) );
  DLY1X1TH U7 ( .A(in[4]), .Y(n30) );
  AOI33X4 U11 ( .A0(n32), .A1(n33), .A2(n23), .B0(n34), .B1(in[5]), .B2(in[4]), 
        .Y(n31) );
  CLKINVX40 U21 ( .A(n31), .Y(n8) );
  CLKINVX40 U22 ( .A(n30), .Y(n32) );
  CLKINVX40 U23 ( .A(in[6]), .Y(n33) );
  AOI21BX4 U24 ( .A0(n25), .A1(n9), .B0N(in[6]), .Y(n34) );
endmodule


module tc_sm_148 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n18, n19, n21, n22, n23, n25, n26, n27,
         n28, n29;

  OAI221XL U4 ( .A0(n18), .A1(n12), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[1])
         );
  OAI221XL U5 ( .A0(n18), .A1(n10), .B0(in[6]), .B1(n22), .C0(n8), .Y(out[2])
         );
  OAI211X1TH U6 ( .A0(in[6]), .A1(n21), .B0(n7), .C0(n8), .Y(out[3]) );
  INVXLTH U8 ( .A(in[6]), .Y(n18) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n21) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U12 ( .A(in[5]), .Y(n19) );
  NAND2BXLTH U13 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  XNOR2XLTH U14 ( .A(n22), .B(n11), .Y(n10) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[2]), .Y(n22) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U18 ( .A(in[1]), .Y(n23) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U20 ( .A0(n9), .A1(n21), .B0(in[6]), .Y(n7) );
  DLY1X1TH U3 ( .A(in[4]), .Y(n25) );
  AOI33X4 U7 ( .A0(n27), .A1(n28), .A2(n19), .B0(n29), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U11 ( .A(n26), .Y(n8) );
  CLKINVX40 U21 ( .A(n25), .Y(n27) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n28) );
  AOI21BX4 U23 ( .A0(n21), .A1(n9), .B0N(in[6]), .Y(n29) );
endmodule


module total_3_test_10 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n60, w5_4_, n4, n5, n6, n7, n42, n43, n44, n49, n50, n51, n52, n53,
         n54, n55, n56;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_151 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_150 sm_tc_2 ( .out(b1), .in({b[4:1], n5}) );
  sm_tc_149 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_148 sm_tc_4 ( .out(in1), .in(in) );
  add_37 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3({c1[6:2], n4, c1[0]}), .in(in1) );
  tc_sm_151 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_150 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_149 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_148 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n51), .CK(clk), .RN(n6), .Q(
        up1[0]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up3[4]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n55), .CK(clk), .RN(n7), .Q(
        h) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n52), .CK(clk), .RN(n6), 
        .Q(up1[3]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n52), .CK(clk), .RN(n6), 
        .Q(n60) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n52), .CK(clk), .RN(n6), 
        .Q(up2[4]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n50), .CK(clk), .RN(n7), 
        .Q(up2[0]) );
  SDFFRQX2TH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n56), .CK(clk), .RN(n6), 
        .Q(up3[1]) );
  SDFFRQX1TH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n53), .CK(clk), .RN(n6), 
        .Q(up1[2]) );
  SDFFRQX2TH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n53), .CK(clk), .RN(n6), 
        .Q(up3[2]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n56), .CK(clk), .RN(n7), 
        .Q(up3[0]) );
  SDFFRQX1 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up2[1]) );
  SDFFRQX1 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n52), .CK(clk), .RN(n6), 
        .Q(up2[2]) );
  BUFX2TH U3 ( .A(c1[1]), .Y(n4) );
  BUFX2TH U4 ( .A(b[0]), .Y(n5) );
  CLKBUFX4TH U5 ( .A(rst), .Y(n6) );
  CLKBUFX1TH U6 ( .A(rst), .Y(n7) );
  SDFFRX4 up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n53), .CK(clk), .RN(n6), 
        .Q(up1[4]) );
  SDFFRX4 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n53), .CK(clk), .RN(n6), 
        .Q(up2[3]) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n55), .CK(clk), .RN(n6), 
        .Q(up1[1]) );
  INVXLTH U39 ( .A(test_se), .Y(n42) );
  INVXLTH U40 ( .A(n42), .Y(n43) );
  INVXLTH U41 ( .A(n42), .Y(n44) );
  DLY1X1TH U42 ( .A(n54), .Y(n49) );
  INVXLTH U43 ( .A(n49), .Y(n50) );
  INVXLTH U44 ( .A(n49), .Y(n51) );
  DLY1X1TH U45 ( .A(n43), .Y(n52) );
  DLY1X1TH U46 ( .A(n44), .Y(n53) );
  INVXLTH U47 ( .A(n43), .Y(n54) );
  INVXLTH U48 ( .A(n49), .Y(n55) );
  INVXLTH U49 ( .A(n49), .Y(n56) );
  DLY1X1TH U50 ( .A(n60), .Y(up3[3]) );
endmodule


module sm_tc_147 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n22, n23, n26, n27, n28;

  INVX6 U2 ( .A(in[4]), .Y(n23) );
  BUFX3 U3 ( .A(n5), .Y(n17) );
  NOR2X6 U4 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2XL U5 ( .A(n22), .B(n8), .Y(n5) );
  CLKBUFX1TH U6 ( .A(out[4]), .Y(out[6]) );
  AOI31X2TH U7 ( .A0(n3), .A1(n4), .A2(n17), .B0(n23), .Y(out[4]) );
  XNOR2X2TH U8 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X2 U9 ( .B0(n23), .B1(n6), .A0N(in[1]), .A1N(n23), .Y(out[1]) );
  INVX2TH U10 ( .A(in[2]), .Y(n22) );
  CLKBUFX1TH U12 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2XLTH U13 ( .B0(n23), .B1(n4), .A0N(in[3]), .A1N(n23), .Y(out[3]) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  AND2X8 U11 ( .A(n8), .B(n22), .Y(n26) );
  CLKINVX40 U15 ( .A(n26), .Y(n7) );
  AOI2B1X4 U16 ( .A1N(n28), .A0(in[1]), .B0(n8), .Y(n27) );
  CLKINVX40 U18 ( .A(n27), .Y(n6) );
  CLKINVX40 U19 ( .A(in[0]), .Y(n28) );
  AO2B2BX4 U20 ( .A0(n23), .A1N(n22), .B0(in[4]), .B1N(n17), .Y(out[2]) );
endmodule


module sm_tc_146 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n22, n23;

  BUFX10 U2 ( .A(in[4]), .Y(n18) );
  XNOR2X2 U3 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2XLTH U4 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  NAND2X1 U5 ( .A(n8), .B(n23), .Y(n7) );
  AO21X4 U6 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X8 U7 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKBUFX2TH U8 ( .A(out[4]), .Y(out[5]) );
  OAI22XLTH U9 ( .A0(n18), .A1(n23), .B0(n22), .B1(n5), .Y(out[2]) );
  CLKBUFX1TH U10 ( .A(out[4]), .Y(out[6]) );
  NOR2BXLTH U11 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2BB2X1TH U12 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U13 ( .A(in[0]), .Y(out[0]) );
  AOI31X4TH U14 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  INVX3TH U15 ( .A(n18), .Y(n22) );
  XNOR2X4 U16 ( .A(n23), .B(n8), .Y(n5) );
  CLKINVX1TH U17 ( .A(in[2]), .Y(n23) );
endmodule


module sm_tc_145 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n20, n21, n22, n23, n27;

  BUFX2 U2 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2XLTH U3 ( .B0(n23), .B1(n4), .A0N(in[3]), .A1N(n23), .Y(out[3]) );
  BUFX10 U4 ( .A(in[1]), .Y(n20) );
  NOR2X3 U5 ( .A(n20), .B(in[0]), .Y(n8) );
  XNOR2X1 U6 ( .A(n7), .B(in[3]), .Y(n4) );
  AO21XLTH U7 ( .A0(in[0]), .A1(n20), .B0(n8), .Y(n6) );
  CLKBUFX1TH U8 ( .A(out[4]), .Y(out[6]) );
  INVX2 U9 ( .A(in[4]), .Y(n23) );
  OAI2BB2X1 U10 ( .B0(n23), .B1(n6), .A0N(n20), .A1N(n23), .Y(out[1]) );
  BUFX2TH U11 ( .A(in[0]), .Y(out[0]) );
  OR2XLTH U12 ( .A(in[4]), .B(n27), .Y(n21) );
  OR2XL U13 ( .A(n23), .B(n5), .Y(n22) );
  CLKNAND2X2TH U14 ( .A(n21), .B(n22), .Y(out[2]) );
  INVX10 U15 ( .A(in[2]), .Y(n27) );
  XNOR2X1TH U16 ( .A(n27), .B(n8), .Y(n5) );
  AOI31X4TH U17 ( .A0(n3), .A1(n4), .A2(n5), .B0(n23), .Y(out[4]) );
  NOR2BXLTH U18 ( .AN(n6), .B(in[0]), .Y(n3) );
  NAND2XLTH U19 ( .A(n8), .B(n27), .Y(n7) );
endmodule


module sm_tc_144 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  AOI31X2 U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  XNOR2X1 U3 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI22X1TH U4 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  NOR2X2TH U5 ( .A(in[1]), .B(in[0]), .Y(n8) );
  NAND2XLTH U6 ( .A(n8), .B(n21), .Y(n7) );
  XNOR2X1TH U7 ( .A(n21), .B(n8), .Y(n5) );
  CLKINVX1TH U8 ( .A(in[2]), .Y(n21) );
  AO21XLTH U9 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKINVX2TH U10 ( .A(in[4]), .Y(n22) );
  INVXLTH U11 ( .A(out[4]), .Y(n18) );
  OAI2BB2X1TH U12 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  INVXLTH U13 ( .A(n18), .Y(out[5]) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2BB2X1TH U15 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  INVXLTH U16 ( .A(n18), .Y(out[6]) );
  CLKBUFX1TH U17 ( .A(in[0]), .Y(out[0]) );
endmodule


module add_36_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_36_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n5), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  NAND2XL U1 ( .A(carry[4]), .B(A[4]), .Y(n2) );
  XOR2XL U2 ( .A(n1), .B(carry[4]), .Y(SUM[4]) );
  NAND2X1 U3 ( .A(carry[4]), .B(B[4]), .Y(n3) );
  NAND3X4 U4 ( .A(n2), .B(n3), .C(n4), .Y(carry[5]) );
  AND2XLTH U6 ( .A(B[0]), .B(A[0]), .Y(n5) );
  CLKXOR2X1TH U7 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2XLTH U8 ( .A(B[4]), .B(A[4]), .Y(n1) );
  AND2X8 U5 ( .A(A[4]), .B(B[4]), .Y(n6) );
  CLKINVX40 U9 ( .A(n6), .Y(n4) );
endmodule


module add_36_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_36_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_36_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [6:2] carry;

  XOR2X2 U12 ( .A(B[4]), .B(carry[4]), .Y(n6) );
  NAND2X2 U13 ( .A(A[4]), .B(carry[4]), .Y(n7) );
  NAND2X2 U14 ( .A(A[4]), .B(B[4]), .Y(n8) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX1 U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  NAND2X1 U1 ( .A(n14), .B(carry[5]), .Y(n12) );
  NAND2X4 U2 ( .A(n10), .B(n11), .Y(n13) );
  NAND2X4 U3 ( .A(n12), .B(n13), .Y(SUM[5]) );
  INVX1 U4 ( .A(n14), .Y(n10) );
  CLKINVX1 U5 ( .A(carry[5]), .Y(n11) );
  XNOR2X1 U6 ( .A(B[5]), .B(A[5]), .Y(n14) );
  NAND3X4 U7 ( .A(n7), .B(n8), .C(n9), .Y(carry[5]) );
  CLKXOR2X2TH U8 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND3X2 U9 ( .A(n3), .B(n4), .C(n5), .Y(carry[6]) );
  NAND2XLTH U10 ( .A(A[5]), .B(B[5]), .Y(n5) );
  CLKXOR2X4TH U11 ( .A(n6), .B(A[4]), .Y(SUM[4]) );
  CLKNAND2X2 U15 ( .A(carry[5]), .B(A[5]), .Y(n3) );
  NAND2XLTH U16 ( .A(carry[5]), .B(B[5]), .Y(n4) );
  AND2XLTH U17 ( .A(B[0]), .B(A[0]), .Y(n1) );
  NAND2X2 U18 ( .A(carry[4]), .B(B[4]), .Y(n9) );
endmodule


module add_36_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_36 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n17, n18, n19, n20, n21;

  add_36_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in2[6:4], n18, n21, in2[1:0]}), 
        .SUM(out3) );
  add_36_DW01_add_1 add_33 ( .A({temp2_6_, n20, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_36_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in3[6:4], n17, in3[2], n19, in3[0]}), .SUM(out2) );
  add_36_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({temp2_6_, n20, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_36_DW01_add_4 add_30 ( .A({in2[6:4], n18, n21, in2[1:0]}), .B({in3[6:4], 
        n17, in3[2], n19, in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_36_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX16 U1 ( .A(temp2_5_), .Y(n20) );
  BUFX4 U2 ( .A(in3[3]), .Y(n17) );
  BUFX4 U3 ( .A(in2[2]), .Y(n21) );
  BUFX4 U4 ( .A(in2[3]), .Y(n18) );
  BUFX8 U5 ( .A(in3[1]), .Y(n19) );
endmodule


module tc_sm_147 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n28, n29, n30, n31, n32, n33;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n33) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n32) );
  XNOR2XLTH U7 ( .A(n32), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(in[4]), .Y(n30) );
  INVXLTH U10 ( .A(in[5]), .Y(n29) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n31) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  OAI33X4TH U13 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n29), .B2(
        n30), .Y(n8) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n28) );
  OAI221XLTH U16 ( .A0(n28), .A1(n12), .B0(in[6]), .B1(n33), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n28), .A1(n10), .B0(in[6]), .B1(n32), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n31), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n31), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n31), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_146 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n22, n25, n27, n28, n29, n30,
         n32, n33, n34, n35;

  CLKBUFX2TH U6 ( .A(in[4]), .Y(n20) );
  NAND3XL U7 ( .A(n21), .B(n22), .C(n8), .Y(out[1]) );
  INVX4 U8 ( .A(n20), .Y(n27) );
  OR2X1TH U9 ( .A(n25), .B(n12), .Y(n21) );
  OR2XLTH U10 ( .A(in[6]), .B(n30), .Y(n22) );
  OAI221X2TH U11 ( .A0(n33), .A1(n10), .B0(in[6]), .B1(n29), .C0(n8), .Y(
        out[2]) );
  OAI211X2TH U12 ( .A0(in[6]), .A1(n28), .B0(n7), .C0(n8), .Y(out[3]) );
  NAND2BX1TH U13 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  CLKINVX1TH U15 ( .A(in[3]), .Y(n28) );
  NOR3X1TH U16 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U17 ( .A(n29), .B(n11), .Y(n10) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U19 ( .A(in[2]), .Y(n29) );
  INVXLTH U20 ( .A(in[1]), .Y(n30) );
  XNOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n12) );
  CLKBUFX1TH U22 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U23 ( .A0(n9), .A1(n28), .B0(in[6]), .Y(n7) );
  INVXLTH U24 ( .A(in[6]), .Y(n25) );
  AOI33X4 U3 ( .A0(n27), .A1(n33), .A2(n34), .B0(n35), .B1(in[5]), .B2(n20), 
        .Y(n32) );
  CLKINVX40 U4 ( .A(n32), .Y(n8) );
  CLKINVX40 U5 ( .A(in[6]), .Y(n33) );
  CLKINVX40 U14 ( .A(in[5]), .Y(n34) );
  AOI21BX4 U25 ( .A0(n28), .A1(n9), .B0N(in[6]), .Y(n35) );
endmodule


module tc_sm_145 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n26, n27,
         n28;

  OAI211X2 U3 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221X2 U5 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1])
         );
  NAND2BX2TH U6 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221X2 U7 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2])
         );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n22) );
  OAI21XLTH U10 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  INVXLTH U11 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U13 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U15 ( .A(in[2]), .Y(n23) );
  CLKBUFX1TH U16 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U17 ( .A(in[6]), .Y(n19) );
  INVX2 U18 ( .A(in[5]), .Y(n20) );
  INVXL U20 ( .A(in[4]), .Y(n21) );
  AOI33X4 U4 ( .A0(n21), .A1(n27), .A2(n20), .B0(n28), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U19 ( .A(n26), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n27) );
  AOI21BX4 U22 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n28) );
endmodule


module tc_sm_144 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n26, n27,
         n28;

  OAI211X1 U3 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221X1 U4 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1])
         );
  NAND2BXL U5 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221X1 U7 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2])
         );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n22) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U11 ( .A(in[4]), .Y(n21) );
  INVXLTH U12 ( .A(in[5]), .Y(n20) );
  INVXLTH U13 ( .A(in[6]), .Y(n19) );
  OAI21XLTH U14 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U16 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U18 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U20 ( .A(in[2]), .Y(n23) );
  AOI33X4 U6 ( .A0(n21), .A1(n27), .A2(n20), .B0(n28), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U8 ( .A(n26), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n27) );
  AOI21BX4 U22 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n28) );
endmodule


module total_3_test_11 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n54, w5_4_, n4, n5, n40, n41, n42, n43, n44, n45, n46, n47, n48, n52,
         n53;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_147 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_146 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_145 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_144 sm_tc_4 ( .out(in1), .in(in) );
  add_36 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_147 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_146 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_145 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_144 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n42), .CK(clk), .RN(n5), .Q(
        up1[0]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n44), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRQX1TH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n43), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n43), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n45), .CK(clk), .RN(n5), .Q(
        h) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up3[3]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n42), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n45), .CK(clk), .RN(n4), 
        .Q(n54) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n44), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n45), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRQXLTH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n44), .CK(clk), .RN(n4), 
        .Q(up1[1]) );
  SDFFRHQX2 up2_reg_4_ ( .D(w7[4]), .SI(n53), .SE(n45), .CK(clk), .RN(n5), .Q(
        up2[4]) );
  SDFFRQX2 up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up1[4]) );
  CLKBUFX4TH U3 ( .A(rst), .Y(n4) );
  CLKBUFX1TH U4 ( .A(rst), .Y(n5) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n44), .CK(clk), .RN(n4), 
        .Q(up1[2]) );
  INVXLTH U37 ( .A(n46), .Y(n40) );
  DLY1X1TH U38 ( .A(n46), .Y(n41) );
  INVXLTH U39 ( .A(n41), .Y(n42) );
  INVXLTH U40 ( .A(n41), .Y(n43) );
  DLY1X1TH U41 ( .A(n40), .Y(n44) );
  DLY1X1TH U42 ( .A(test_se), .Y(n45) );
  INVXLTH U43 ( .A(test_se), .Y(n46) );
  INVXLTH U44 ( .A(n41), .Y(n47) );
  INVXLTH U45 ( .A(n41), .Y(n48) );
  DLY1X1TH U46 ( .A(n54), .Y(up2[3]) );
  INVXLTH U47 ( .A(up2[3]), .Y(n52) );
  INVXLTH U48 ( .A(n52), .Y(n53) );
endmodule


module sm_tc_143 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n17, n19, n20, n24, n25, n28, n29, n30;

  NAND2X2TH U4 ( .A(n17), .B(n28), .Y(n20) );
  CLKNAND2X4TH U5 ( .A(n19), .B(n20), .Y(n5) );
  AOI31X2TH U6 ( .A0(n3), .A1(n4), .A2(n5), .B0(n24), .Y(out[4]) );
  AO21X1TH U7 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2X4 U9 ( .B0(n24), .B1(n6), .A0N(in[1]), .A1N(n24), .Y(out[1]) );
  NAND2XLTH U10 ( .A(n25), .B(n8), .Y(n19) );
  INVXLTH U11 ( .A(n25), .Y(n17) );
  INVX2TH U13 ( .A(in[2]), .Y(n25) );
  OAI2BB2X1 U14 ( .B0(n24), .B1(n4), .A0N(in[3]), .A1N(n24), .Y(out[3]) );
  INVX4TH U16 ( .A(in[4]), .Y(n24) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX1TH U18 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U19 ( .AN(n6), .B(in[0]), .Y(n3) );
  BUFX2TH U20 ( .A(in[0]), .Y(out[0]) );
  OR2X8 U2 ( .A(in[1]), .B(in[0]), .Y(n28) );
  CLKINVX40 U3 ( .A(n28), .Y(n8) );
  XOR2X1 U8 ( .A(n29), .B(in[3]), .Y(n4) );
  CLKAND2X12 U12 ( .A(n8), .B(n25), .Y(n29) );
  AO2B2BX4 U15 ( .A0(n24), .A1N(n25), .B0(n30), .B1N(n5), .Y(out[2]) );
  CLKINVX40 U21 ( .A(n24), .Y(n30) );
endmodule


module sm_tc_142 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n23, n25, n26, n27, n31, n32, n35;

  BUFX10 U2 ( .A(in[4]), .Y(n23) );
  INVX6 U3 ( .A(n23), .Y(n31) );
  NOR2X3 U4 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKNAND2X2 U5 ( .A(n7), .B(in[3]), .Y(n26) );
  OAI2BB2XL U6 ( .B0(n31), .B1(n4), .A0N(in[3]), .A1N(n31), .Y(out[3]) );
  OAI22X1 U7 ( .A0(n23), .A1(n32), .B0(n31), .B1(n5), .Y(out[2]) );
  CLKNAND2X2TH U9 ( .A(n35), .B(n25), .Y(n27) );
  INVXLTH U10 ( .A(in[3]), .Y(n25) );
  OAI2BB2X2TH U11 ( .B0(n31), .B1(n6), .A0N(in[1]), .A1N(n31), .Y(out[1]) );
  NAND2X4TH U12 ( .A(n26), .B(n27), .Y(n4) );
  INVX1TH U13 ( .A(in[2]), .Y(n32) );
  CLKBUFX1TH U15 ( .A(in[0]), .Y(out[0]) );
  AOI31X4 U16 ( .A0(n3), .A1(n4), .A2(n5), .B0(n31), .Y(out[4]) );
  NOR2BXLTH U18 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U19 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U20 ( .A(out[4]), .Y(out[6]) );
  AO21XLTH U21 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  XOR2X1 U8 ( .A(in[2]), .B(n8), .Y(n5) );
  AND2X8 U14 ( .A(n8), .B(n32), .Y(n35) );
  CLKINVX40 U17 ( .A(n35), .Y(n7) );
endmodule


module sm_tc_141 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n23, n26, n27;

  NOR2X2TH U4 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX6TH U5 ( .A(in[4]), .Y(n23) );
  XNOR2X4 U6 ( .A(n7), .B(in[3]), .Y(n4) );
  XNOR2X1 U7 ( .A(n22), .B(n8), .Y(n5) );
  INVX1TH U8 ( .A(in[2]), .Y(n22) );
  CLKBUFX1TH U9 ( .A(out[4]), .Y(out[6]) );
  AO21X1 U10 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2XLTH U11 ( .B0(n23), .B1(n4), .A0N(in[3]), .A1N(n23), .Y(out[3]) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[5]) );
  AOI31X4TH U14 ( .A0(n3), .A1(n4), .A2(n5), .B0(n23), .Y(out[4]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  BUFX2TH U16 ( .A(in[0]), .Y(out[0]) );
  AND2X8 U2 ( .A(n8), .B(n22), .Y(n26) );
  CLKINVX40 U3 ( .A(n26), .Y(n7) );
  AO2B2X4 U12 ( .B0(in[1]), .B1(n23), .A0(in[4]), .A1N(n6), .Y(out[1]) );
  OAI2B2X2 U17 ( .A1N(n27), .A0(n5), .B0(in[4]), .B1(n22), .Y(out[2]) );
  CLKINVX40 U18 ( .A(n23), .Y(n27) );
endmodule


module sm_tc_140 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  OAI2BB2X2 U2 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  OAI22X1TH U3 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  INVX1TH U4 ( .A(out[4]), .Y(n18) );
  OAI2BB2X1TH U5 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U6 ( .A(in[0]), .Y(out[0]) );
  CLKNAND2X2TH U7 ( .A(n8), .B(n21), .Y(n7) );
  CLKINVX2TH U8 ( .A(in[4]), .Y(n22) );
  NOR2X3TH U9 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X1TH U10 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n21) );
  XNOR2X1TH U12 ( .A(n21), .B(n8), .Y(n5) );
  AOI31X2TH U13 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U15 ( .A(n18), .Y(out[5]) );
  INVXLTH U16 ( .A(n18), .Y(out[6]) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_35_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_35_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [6:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3XLTH U1 ( .A(carry[3]), .B(A[3]), .C(B[3]), .Y(SUM[3]) );
  CLKNAND2X4TH U2 ( .A(carry[3]), .B(A[3]), .Y(n3) );
  CLKNAND2X4TH U3 ( .A(carry[3]), .B(B[3]), .Y(n4) );
  NAND2X2 U4 ( .A(A[3]), .B(B[3]), .Y(n5) );
  NAND3X8 U5 ( .A(n3), .B(n4), .C(n5), .Y(carry[4]) );
  CLKNAND2X12 U6 ( .A(n8), .B(n9), .Y(SUM[6]) );
  NAND2X4 U7 ( .A(n6), .B(n7), .Y(n9) );
  XNOR2X4 U8 ( .A(B[6]), .B(A[6]), .Y(n10) );
  CLKNAND2X2 U9 ( .A(n10), .B(carry[6]), .Y(n8) );
  CLKINVX4 U10 ( .A(n10), .Y(n6) );
  CLKXOR2X1TH U11 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  INVXLTH U12 ( .A(carry[6]), .Y(n7) );
  AND2XLTH U13 ( .A(B[0]), .B(A[0]), .Y(n2) );
endmodule


module add_35_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_35_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX4TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_35_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [6:2] carry;

  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  NAND2X2 U1 ( .A(n8), .B(n9), .Y(SUM[4]) );
  INVX12 U2 ( .A(n2), .Y(n6) );
  CLKNAND2X4 U3 ( .A(n2), .B(n7), .Y(n8) );
  XOR2X8 U4 ( .A(A[4]), .B(B[4]), .Y(n2) );
  NAND3X2 U5 ( .A(n3), .B(n4), .C(n5), .Y(carry[5]) );
  CLKNAND2X2 U6 ( .A(n6), .B(carry[4]), .Y(n9) );
  CLKXOR2X1TH U7 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  INVXLTH U8 ( .A(carry[4]), .Y(n7) );
  NAND2XLTH U9 ( .A(B[4]), .B(A[4]), .Y(n5) );
  NAND2XLTH U10 ( .A(carry[4]), .B(B[4]), .Y(n3) );
  NAND2XLTH U11 ( .A(carry[4]), .B(A[4]), .Y(n4) );
  AND2XLTH U12 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_35_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_35 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31;

  add_35_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n31, n30, 
        temp1_1_, temp1_0_}), .B({in2[6:4], n24, in2[2:0]}), .SUM(out3) );
  add_35_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, n23, temp2_3_, n26, 
        temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_35_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n31, n30, 
        temp1_1_, temp1_0_}), .B({in3[6:4], n29, n22, n25, in3[0]}), .SUM(out2) );
  add_35_DW01_add_3 add_31 ( .A({temp1_6_, n21, temp1_4_, n31, n30, n28, 
        temp1_0_}), .B({temp2_6_, temp2_5_, n23, temp2_3_, n26, temp2_1_, 
        temp2_0_}), .SUM(out) );
  add_35_DW01_add_4 add_30 ( .A({in2[6:4], n24, in2[2:0]}), .B({in3[6:4], n29, 
        n22, in3[1:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}) );
  add_35_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX2TH U1 ( .A(temp1_5_), .Y(n21) );
  BUFX4 U2 ( .A(in3[2]), .Y(n22) );
  BUFX2 U3 ( .A(temp2_4_), .Y(n23) );
  CLKBUFX1TH U4 ( .A(temp2_2_), .Y(n26) );
  BUFX2 U5 ( .A(in2[3]), .Y(n24) );
  BUFX2TH U6 ( .A(in3[1]), .Y(n25) );
  INVXLTH U13 ( .A(temp1_1_), .Y(n27) );
  INVXLTH U14 ( .A(n27), .Y(n28) );
  CLKBUFX1TH U15 ( .A(in3[3]), .Y(n29) );
  CLKBUFX40 U16 ( .A(temp1_2_), .Y(n30) );
  CLKBUFX40 U17 ( .A(temp1_3_), .Y(n31) );
endmodule


module tc_sm_143 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n27, n28, n29, n30, n31, n32;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n31) );
  XNOR2XLTH U7 ( .A(n31), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n28), .B2(
        n29), .Y(n8) );
  INVXLTH U10 ( .A(in[5]), .Y(n28) );
  INVXLTH U11 ( .A(in[4]), .Y(n29) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n30) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n27) );
  OAI221XLTH U16 ( .A0(n27), .A1(n12), .B0(in[6]), .B1(n32), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n27), .A1(n10), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n30), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n30), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n30), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_142 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n17, n18, n19, n22, n25, n26, n27, n29,
         n30, n31, n32, n33, n34, n35, n36;

  NOR2X2 U3 ( .A(n32), .B(n10), .Y(n17) );
  NOR2XL U4 ( .A(in[6]), .B(n26), .Y(n18) );
  CLKINVX1 U5 ( .A(n8), .Y(n19) );
  OR3X4 U6 ( .A(n17), .B(n18), .C(n19), .Y(out[2]) );
  XNOR2X1 U7 ( .A(n26), .B(n11), .Y(n10) );
  CLKINVX2TH U8 ( .A(in[2]), .Y(n26) );
  INVXLTH U10 ( .A(in[6]), .Y(n22) );
  OAI221X2TH U13 ( .A0(n22), .A1(n12), .B0(in[6]), .B1(n27), .C0(n8), .Y(
        out[1]) );
  CLKINVX1TH U15 ( .A(in[3]), .Y(n25) );
  NOR3X1TH U16 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U18 ( .A(in[1]), .Y(n27) );
  XNOR2XLTH U19 ( .A(n29), .B(in[1]), .Y(n12) );
  NOR2XLTH U20 ( .A(n29), .B(in[1]), .Y(n11) );
  OAI21XLTH U21 ( .A0(n9), .A1(n25), .B0(in[6]), .Y(n7) );
  INVXLTH U9 ( .A(n36), .Y(n29) );
  OAI2B11X4 U11 ( .A1N(n32), .A0(n25), .B0(n7), .C0(n8), .Y(out[3]) );
  AOI33X4 U12 ( .A0(n31), .A1(n32), .A2(n33), .B0(n34), .B1(in[5]), .B2(in[4]), 
        .Y(n30) );
  CLKINVX40 U14 ( .A(n30), .Y(n8) );
  CLKINVX40 U22 ( .A(in[4]), .Y(n31) );
  CLKINVX40 U23 ( .A(in[6]), .Y(n32) );
  CLKINVX40 U24 ( .A(in[5]), .Y(n33) );
  AOI21BX4 U25 ( .A0(n25), .A1(n9), .B0N(in[6]), .Y(n34) );
  AND2X8 U26 ( .A(n36), .B(n8), .Y(n35) );
  CLKINVX40 U27 ( .A(n35), .Y(out[0]) );
  CLKINVX40 U28 ( .A(in[0]), .Y(n36) );
endmodule


module tc_sm_141 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n22, n23, n24, n26, n27, n28,
         n29, n30, n31;

  OAI211XL U3 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221XL U5 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2])
         );
  OAI221XL U6 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1])
         );
  NOR3X1TH U7 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n22) );
  INVXLTH U9 ( .A(in[6]), .Y(n19) );
  NAND2BXLTH U10 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  CLKBUFX1TH U11 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U12 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  XNOR2XLTH U13 ( .A(n23), .B(n11), .Y(n10) );
  INVX2 U14 ( .A(in[5]), .Y(n20) );
  INVXLTH U15 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U18 ( .A(in[2]), .Y(n23) );
  DLY1X1TH U4 ( .A(in[4]), .Y(n26) );
  AOI33X4 U19 ( .A0(n28), .A1(n29), .A2(n20), .B0(n31), .B1(n30), .B2(in[4]), 
        .Y(n27) );
  CLKINVX40 U20 ( .A(n27), .Y(n8) );
  CLKINVX40 U21 ( .A(n26), .Y(n28) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n29) );
  CLKINVX40 U23 ( .A(n20), .Y(n30) );
  AOI21BX4 U24 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n31) );
endmodule


module tc_sm_140 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n24, n25, n27, n28, n29, n30;

  OAI221XL U3 ( .A0(n27), .A1(n10), .B0(in[6]), .B1(n30), .C0(n6), .Y(out[1])
         );
  CLKAND2X3TH U4 ( .A(n25), .B(n24), .Y(n6) );
  NAND2XLTH U5 ( .A(in[6]), .B(n11), .Y(n25) );
  OAI2B11X2TH U6 ( .A1N(n7), .A0(in[3]), .B0(in[5]), .C0(in[4]), .Y(n11) );
  OAI221XLTH U7 ( .A0(n27), .A1(n8), .B0(in[6]), .B1(n29), .C0(n6), .Y(out[2])
         );
  OAI211XLTH U8 ( .A0(in[6]), .A1(n28), .B0(n5), .C0(n6), .Y(out[3]) );
  NAND2BXLTH U9 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  OAI21BXLTH U10 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n24) );
  INVXLTH U11 ( .A(in[6]), .Y(n27) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  INVXLTH U13 ( .A(in[2]), .Y(n29) );
  XOR2XLTH U14 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n9) );
  XOR2XLTH U16 ( .A(in[0]), .B(n30), .Y(n10) );
  INVXLTH U17 ( .A(in[1]), .Y(n30) );
  OAI21XLTH U18 ( .A0(n7), .A1(n28), .B0(in[6]), .Y(n5) );
  INVXLTH U19 ( .A(in[3]), .Y(n28) );
  CLKBUFX1TH U20 ( .A(in[6]), .Y(out[4]) );
endmodule


module total_3_test_12 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n4, n39, n40, n41, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_143 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_142 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_141 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_140 sm_tc_4 ( .out(in1), .in(in) );
  add_35 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_143 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_142 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_141 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_140 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n52), .CK(clk), .RN(n4), .Q(
        h) );
  SDFFRHQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up1[4]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRQX1TH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n49), .CK(clk), .RN(rst), 
        .Q(up1[1]) );
  SDFFRHQX1TH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  SDFFRHQX1TH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRHQX1TH up2_reg_1_ ( .D(w7[1]), .SI(n55), .SE(n53), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n50), .CK(clk), .RN(n4), .Q(
        up1[0]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRQX2TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRHQX1TH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up2[3]) );
  SDFFRQX2 up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up2[4]) );
  SDFFRHQX2 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up1[2]) );
  CLKBUFX4TH U3 ( .A(rst), .Y(n4) );
  SDFFRX4 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n53), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRX4 up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up3[3]) );
  INVXLTH U36 ( .A(test_se), .Y(n39) );
  INVXLTH U37 ( .A(n39), .Y(n40) );
  INVXLTH U38 ( .A(n39), .Y(n41) );
  DLY1X1TH U39 ( .A(n51), .Y(n46) );
  INVXLTH U40 ( .A(n46), .Y(n47) );
  INVXLTH U41 ( .A(n46), .Y(n48) );
  DLY1X1TH U42 ( .A(n40), .Y(n49) );
  DLY1X1TH U43 ( .A(n41), .Y(n50) );
  INVXLTH U44 ( .A(n40), .Y(n51) );
  INVXLTH U45 ( .A(n46), .Y(n52) );
  INVXLTH U46 ( .A(n46), .Y(n53) );
  INVXLTH U47 ( .A(up2[0]), .Y(n54) );
  INVXLTH U48 ( .A(n54), .Y(n55) );
endmodule


module sm_tc_139 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n23, n27, n28, n31, n32;

  BUFX2 U2 ( .A(in[4]), .Y(n23) );
  BUFX2TH U3 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U4 ( .A(out[4]), .Y(out[6]) );
  NOR2X2 U5 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X2TH U6 ( .A(n27), .B(n8), .Y(n5) );
  OAI2BB2X4TH U7 ( .B0(n32), .B1(n6), .A0N(in[1]), .A1N(n32), .Y(out[1]) );
  AOI31X2TH U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n32), .Y(out[4]) );
  XNOR2X4 U9 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX3TH U10 ( .A(n23), .Y(n28) );
  INVX1TH U11 ( .A(in[2]), .Y(n27) );
  OAI2BB2XLTH U12 ( .B0(n32), .B1(n4), .A0N(in[3]), .A1N(n32), .Y(out[3]) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  AO21X2 U15 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI22XLTH U16 ( .A0(n23), .A1(n27), .B0(n32), .B1(n5), .Y(out[2]) );
  NAND2XLTH U17 ( .A(n8), .B(n27), .Y(n7) );
  CLKINVX40 U18 ( .A(n28), .Y(n31) );
  CLKINVX40 U19 ( .A(n31), .Y(n32) );
endmodule


module sm_tc_138 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n20, n21, n24, n25, n26, n27, n28;

  OAI2BB2X2 U5 ( .B0(n20), .B1(n6), .A0N(in[1]), .A1N(n20), .Y(out[1]) );
  AO21X2 U2 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  BUFX2 U3 ( .A(in[0]), .Y(out[0]) );
  NOR2X4 U4 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKBUFX1TH U6 ( .A(out[4]), .Y(out[6]) );
  INVX4TH U7 ( .A(in[4]), .Y(n20) );
  INVX2TH U10 ( .A(in[2]), .Y(n21) );
  OAI22X2TH U11 ( .A0(n26), .A1(n21), .B0(n20), .B1(n5), .Y(out[2]) );
  AOI31X2TH U14 ( .A0(n3), .A1(n4), .A2(n27), .B0(n20), .Y(out[4]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  OAI2B2X2 U8 ( .A1N(in[3]), .A0(n24), .B0(n20), .B1(n4), .Y(out[3]) );
  CLKINVX40 U9 ( .A(n20), .Y(n24) );
  XOR2X1 U12 ( .A(n25), .B(in[3]), .Y(n4) );
  CLKAND2X12 U13 ( .A(n8), .B(n21), .Y(n25) );
  CLKINVX40 U17 ( .A(n20), .Y(n26) );
  XOR2X1 U18 ( .A(n21), .B(n28), .Y(n27) );
  XOR2X1 U19 ( .A(n21), .B(n28), .Y(n5) );
  CLKINVX40 U20 ( .A(n8), .Y(n28) );
endmodule


module sm_tc_137 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n23, n24, n28, n29, n32, n33;

  BUFX5 U2 ( .A(in[0]), .Y(n22) );
  OAI2BB2X1TH U4 ( .B0(n29), .B1(n6), .A0N(n24), .A1N(n29), .Y(out[1]) );
  OAI22X4 U5 ( .A0(n23), .A1(n28), .B0(n29), .B1(n5), .Y(out[2]) );
  AOI31X2 U6 ( .A0(n3), .A1(n4), .A2(n5), .B0(n29), .Y(out[4]) );
  OAI2BB2X2TH U7 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  INVX8 U8 ( .A(n23), .Y(n29) );
  BUFX4 U9 ( .A(in[4]), .Y(n23) );
  XNOR2X2 U10 ( .A(n28), .B(n8), .Y(n5) );
  XNOR2X2TH U11 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX2TH U12 ( .A(in[1]), .Y(n24) );
  CLKBUFX1TH U13 ( .A(n22), .Y(out[0]) );
  INVX1TH U14 ( .A(in[2]), .Y(n28) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[6]) );
  NOR2BXLTH U16 ( .AN(n6), .B(n22), .Y(n3) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[5]) );
  NAND2XLTH U18 ( .A(n8), .B(n28), .Y(n7) );
  OR2X8 U3 ( .A(n24), .B(n22), .Y(n32) );
  CLKINVX40 U19 ( .A(n32), .Y(n8) );
  AOI21BX4 U20 ( .A0(n22), .A1(n24), .B0N(n32), .Y(n33) );
  CLKINVX40 U21 ( .A(n33), .Y(n6) );
endmodule


module sm_tc_136 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n20, n21;

  OAI2BB2X2 U5 ( .B0(n21), .B1(n6), .A0N(in[1]), .A1N(n21), .Y(out[1]) );
  CLKBUFX1TH U2 ( .A(in[0]), .Y(out[0]) );
  NOR2X2TH U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  NAND2X1TH U4 ( .A(n8), .B(n20), .Y(n7) );
  OAI2BB2X2TH U6 ( .B0(n21), .B1(n4), .A0N(in[3]), .A1N(n21), .Y(out[3]) );
  AOI31X4TH U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n21), .Y(out[6]) );
  OAI22X1TH U8 ( .A0(in[4]), .A1(n20), .B0(n21), .B1(n5), .Y(out[2]) );
  CLKINVX2TH U9 ( .A(in[4]), .Y(n21) );
  NOR2BXLTH U10 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n20) );
  CLKBUFX1TH U12 ( .A(out[6]), .Y(out[5]) );
  CLKBUFX1TH U13 ( .A(out[6]), .Y(out[4]) );
  XNOR2X1TH U14 ( .A(n20), .B(n8), .Y(n5) );
  XNOR2X1TH U15 ( .A(n7), .B(in[3]), .Y(n4) );
  AO21XLTH U16 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_34_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n8, n1, n2, n3, n4, n5, n6;
  wire   [6:2] carry;

  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n8) );
  ADDFX2TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  NAND2XL U2 ( .A(carry[2]), .B(B[2]), .Y(n4) );
  NAND3X2TH U3 ( .A(n3), .B(n4), .C(n5), .Y(carry[3]) );
  XOR2XLTH U4 ( .A(B[2]), .B(A[2]), .Y(n2) );
  CLKXOR2X1TH U5 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2XLTH U6 ( .A(A[2]), .B(B[2]), .Y(n5) );
  NAND2XLTH U7 ( .A(carry[2]), .B(A[2]), .Y(n3) );
  XOR2X1TH U8 ( .A(n2), .B(carry[2]), .Y(SUM[2]) );
  CLKINVX40 U9 ( .A(n8), .Y(n6) );
  CLKINVX40 U10 ( .A(n6), .Y(SUM[6]) );
endmodule


module add_34_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_34_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_34_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_34_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_34_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_34 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n17, n18, n19, n20, n21, n22;

  add_34_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in2[6:3], n19, in2[1:0]}), .SUM(
        out3) );
  add_34_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, n21, temp2_3_, n20, 
        temp2_1_, n22}), .B(in), .SUM(out1) );
  add_34_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in3[6:3], n18, n17, in3[0]}), 
        .SUM(out2) );
  add_34_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, n21, temp2_3_, 
        n20, temp2_1_, n22}), .SUM(out) );
  add_34_DW01_add_4 add_30 ( .A({in2[6:3], n19, in2[1:0]}), .B({in3[6:3], n18, 
        n17, in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_34_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX6 U1 ( .A(in3[1]), .Y(n17) );
  BUFX2TH U2 ( .A(in3[2]), .Y(n18) );
  CLKBUFX16 U3 ( .A(in2[2]), .Y(n19) );
  CLKBUFX40 U4 ( .A(temp2_2_), .Y(n20) );
  CLKBUFX40 U5 ( .A(temp2_4_), .Y(n21) );
  CLKBUFX40 U6 ( .A(temp2_0_), .Y(n22) );
endmodule


module tc_sm_139 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U10 ( .A(in[4]), .Y(n28) );
  INVXLTH U11 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI2BB1XLTH U19 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI211XLTH U20 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
endmodule


module tc_sm_138 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n19, n20, n21, n22, n24, n25,
         n26, n27, n28, n29;

  NAND3XL U3 ( .A(n19), .B(n20), .C(n22), .Y(out[2]) );
  NAND2XLTH U4 ( .A(n18), .B(n22), .Y(out[3]) );
  OAI221X1TH U5 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n22), .Y(
        out[1]) );
  INVXLTH U6 ( .A(in[6]), .Y(n24) );
  CLKINVX20 U7 ( .A(n21), .Y(n22) );
  OA21XL U8 ( .A0(in[6]), .A1(n27), .B0(n7), .Y(n18) );
  OR2X1 U9 ( .A(n24), .B(n10), .Y(n19) );
  OR2XLTH U10 ( .A(in[6]), .B(n28), .Y(n20) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n27) );
  OAI2BB1X4 U12 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U14 ( .A(in[5]), .Y(n25) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U16 ( .A(n28), .B(n11), .Y(n10) );
  OAI21XLTH U17 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  INVX6 U18 ( .A(n8), .Y(n21) );
  NOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U20 ( .A(in[2]), .Y(n28) );
  INVXLTH U21 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U22 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U23 ( .AN(in[0]), .B(n22), .Y(out[0]) );
  OAI33X4 U24 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXL U25 ( .A(in[4]), .Y(n26) );
endmodule


module tc_sm_137 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n22, n23, n24, n26, n27, n28,
         n29, n30;

  OAI211X2TH U3 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  NAND2BX1TH U5 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221X2TH U6 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1]) );
  OAI221X2TH U7 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2]) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n22) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U10 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U12 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  XNOR2XLTH U13 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U15 ( .A(in[2]), .Y(n23) );
  CLKBUFX1TH U16 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U17 ( .A(in[6]), .Y(n19) );
  INVXL U19 ( .A(in[5]), .Y(n20) );
  INVXLTH U4 ( .A(n28), .Y(n26) );
  AOI33X4 U18 ( .A0(n28), .A1(n29), .A2(n20), .B0(n30), .B1(in[5]), .B2(n26), 
        .Y(n27) );
  CLKINVX40 U20 ( .A(n27), .Y(n8) );
  CLKINVX40 U21 ( .A(in[4]), .Y(n28) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n29) );
  AOI21BX4 U23 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n30) );
endmodule


module tc_sm_136 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n23, n24, n25, n26, n28, n29, n30, n31,
         n32;

  INVX4 U3 ( .A(n23), .Y(n8) );
  INVXL U4 ( .A(in[6]), .Y(n25) );
  INVXLTH U5 ( .A(in[4]), .Y(n24) );
  AOI33X4 U6 ( .A0(n24), .A1(n25), .A2(n30), .B0(n26), .B1(in[5]), .B2(in[4]), 
        .Y(n23) );
  AOI21BX2 U7 ( .A0(n31), .A1(n9), .B0N(in[6]), .Y(n26) );
  OAI211XLTH U8 ( .A0(in[6]), .A1(n31), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221XLTH U9 ( .A0(n29), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(out[2]) );
  OAI221XLTH U10 ( .A0(n29), .A1(n12), .B0(in[6]), .B1(n32), .C0(n8), .Y(
        out[1]) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n31) );
  INVXLTH U12 ( .A(in[6]), .Y(n29) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U14 ( .A(n28), .B(n11), .Y(n10) );
  OAI21XLTH U15 ( .A0(n9), .A1(n31), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U16 ( .A(in[6]), .Y(out[4]) );
  INVX2 U17 ( .A(in[5]), .Y(n30) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U19 ( .A(in[2]), .Y(n28) );
  INVXLTH U20 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U22 ( .AN(in[0]), .B(n8), .Y(out[0]) );
endmodule


module total_3_test_13 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n5, n6, n41, n42, n43, n44, n45, n46, n47, n48, n49;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_139 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_138 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_137 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_136 sm_tc_4 ( .out(in1), .in(in) );
  add_34 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_139 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_138 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_137 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_136 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n44), .CK(clk), .RN(n5), 
        .Q(up3[3]) );
  SDFFRQX4TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n43), .CK(clk), .RN(n6), 
        .Q(up2[1]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n45), .CK(clk), .RN(n5), .Q(
        up1[0]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n44), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n45), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  SDFFRQX1TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up3[4]) );
  SDFFRQX2 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n45), .CK(clk), .RN(n5), 
        .Q(up1[2]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n43), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRQX2 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n6) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n5) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up1[1]) );
  SDFFRX4 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up2[2]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up1[3]) );
  SDFFRX4 h_reg ( .D(w5_4_), .SI(test_si), .SE(n45), .CK(clk), .RN(n6), .Q(h)
         );
  INVXLTH U37 ( .A(n47), .Y(n41) );
  DLY1X1TH U38 ( .A(n47), .Y(n42) );
  INVXLTH U39 ( .A(n42), .Y(n43) );
  INVXLTH U40 ( .A(n42), .Y(n44) );
  DLY1X1TH U41 ( .A(n41), .Y(n45) );
  DLY1X1TH U42 ( .A(test_se), .Y(n46) );
  INVXLTH U43 ( .A(test_se), .Y(n47) );
  INVXLTH U44 ( .A(n42), .Y(n48) );
  INVXLTH U45 ( .A(n42), .Y(n49) );
endmodule


module sm_tc_135 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n29, n33, n34, n37, n38;

  BUFX2 U2 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X4 U4 ( .B0(n33), .B1(n6), .A0N(n37), .A1N(n33), .Y(out[1]) );
  BUFX6 U5 ( .A(in[4]), .Y(n29) );
  NOR2X6 U6 ( .A(n37), .B(in[0]), .Y(n8) );
  INVX2TH U8 ( .A(in[2]), .Y(n34) );
  XNOR2X2TH U9 ( .A(n34), .B(n8), .Y(n5) );
  AO21X2TH U10 ( .A0(in[0]), .A1(n37), .B0(n8), .Y(n6) );
  INVX2TH U11 ( .A(n29), .Y(n33) );
  OAI2BB2X1TH U12 ( .B0(n33), .B1(n4), .A0N(in[3]), .A1N(n33), .Y(out[3]) );
  AOI31X2TH U13 ( .A0(n3), .A1(n4), .A2(n5), .B0(n33), .Y(out[4]) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[6]) );
  OAI22X1TH U15 ( .A0(n29), .A1(n34), .B0(n33), .B1(n5), .Y(out[2]) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX40 U3 ( .A(in[1]), .Y(n37) );
  XOR2X1 U7 ( .A(n38), .B(in[3]), .Y(n4) );
  CLKAND2X12 U18 ( .A(n8), .B(n34), .Y(n38) );
endmodule


module sm_tc_134 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n19, n20, n21, n22, n26, n27, n30, n31;

  XNOR2X1 U2 ( .A(n7), .B(n31), .Y(n4) );
  NAND3X4 U3 ( .A(n3), .B(n4), .C(n5), .Y(n22) );
  NAND2XLTH U6 ( .A(n27), .B(n8), .Y(n20) );
  NAND2X2 U7 ( .A(n18), .B(n19), .Y(n21) );
  NAND2X4 U8 ( .A(n20), .B(n21), .Y(n5) );
  INVXLTH U9 ( .A(n27), .Y(n18) );
  INVXLTH U10 ( .A(n8), .Y(n19) );
  INVX4 U11 ( .A(in[2]), .Y(n27) );
  NOR2X6 U12 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI22X2 U13 ( .A0(in[4]), .A1(n27), .B0(n26), .B1(n5), .Y(out[2]) );
  AND2X1TH U14 ( .A(n22), .B(in[4]), .Y(out[4]) );
  INVX2 U15 ( .A(in[4]), .Y(n26) );
  BUFX2TH U16 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U18 ( .A(out[4]), .Y(out[6]) );
  AO21XLTH U19 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2BXLTH U20 ( .AN(n6), .B(in[0]), .Y(n3) );
  NAND2XLTH U21 ( .A(n8), .B(n27), .Y(n7) );
  AO2B2X4 U4 ( .B0(in[1]), .B1(n26), .A0(in[4]), .A1N(n6), .Y(out[1]) );
  OAI2B2X2 U5 ( .A1N(n26), .A0(n30), .B0(n26), .B1(n4), .Y(out[3]) );
  CLKINVX40 U22 ( .A(n31), .Y(n30) );
  CLKBUFX40 U23 ( .A(in[3]), .Y(n31) );
endmodule


module sm_tc_133 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n37, n3, n4, n5, n6, n7, n8, n29, n30, n33, n35, n36;

  XNOR2X4 U3 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX10 U4 ( .A(n36), .Y(n30) );
  BUFX10 U5 ( .A(in[0]), .Y(out[0]) );
  NOR2X8 U6 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI2BB2X2 U7 ( .B0(n30), .B1(n6), .A0N(in[1]), .A1N(n30), .Y(out[1]) );
  AOI31X2 U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n30), .Y(n37) );
  XNOR2X4 U10 ( .A(n29), .B(n8), .Y(n5) );
  INVX2 U11 ( .A(in[2]), .Y(n29) );
  OAI2BB2X1TH U12 ( .B0(n30), .B1(n4), .A0N(in[3]), .A1N(n30), .Y(out[3]) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[6]) );
  AO21X2 U15 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2BXLTH U16 ( .AN(n6), .B(out[0]), .Y(n3) );
  OAI2BB2X2 U2 ( .B0(n30), .B1(n5), .A0N(n30), .A1N(in[2]), .Y(out[2]) );
  CLKINVX40 U9 ( .A(n37), .Y(n33) );
  CLKINVX40 U17 ( .A(n33), .Y(out[4]) );
  AND2X8 U18 ( .A(n8), .B(n29), .Y(n35) );
  CLKINVX40 U19 ( .A(n35), .Y(n7) );
  CLKBUFX40 U20 ( .A(in[4]), .Y(n36) );
endmodule


module sm_tc_132 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n19, n22, n23;

  OAI2BB2X2 U5 ( .B0(n23), .B1(n6), .A0N(in[1]), .A1N(n23), .Y(out[1]) );
  AND3X2 U2 ( .A(n3), .B(n4), .C(n5), .Y(n17) );
  NOR2X2 U3 ( .A(n17), .B(n23), .Y(out[4]) );
  XNOR2X1TH U4 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX2TH U6 ( .A(in[0]), .Y(out[0]) );
  CLKINVX1TH U7 ( .A(in[2]), .Y(n22) );
  OAI22X1TH U8 ( .A0(in[4]), .A1(n22), .B0(n23), .B1(n5), .Y(out[2]) );
  NAND2XLTH U9 ( .A(n8), .B(n22), .Y(n7) );
  NOR2X6 U10 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX2TH U11 ( .A(in[4]), .Y(n23) );
  INVXLTH U12 ( .A(n19), .Y(out[6]) );
  XNOR2X1TH U13 ( .A(n22), .B(n8), .Y(n5) );
  INVXLTH U14 ( .A(out[4]), .Y(n19) );
  INVXLTH U15 ( .A(n19), .Y(out[5]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2BB2X1TH U17 ( .B0(n23), .B1(n4), .A0N(in[3]), .A1N(n23), .Y(out[3]) );
  AO21XLTH U18 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_33_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1TH U1_1 ( .A(B[1]), .B(A[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX4TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  NAND3X2 U1 ( .A(n3), .B(n4), .C(n5), .Y(carry[3]) );
  NAND2XL U2 ( .A(carry[2]), .B(B[2]), .Y(n5) );
  CLKXOR2X4 U3 ( .A(n6), .B(carry[6]), .Y(SUM[6]) );
  CLKAND2X2TH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XLTH U5 ( .A(B[6]), .B(A[6]), .Y(n6) );
  CLKXOR2X1TH U6 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2XLTH U7 ( .A(B[2]), .B(carry[2]), .Y(n2) );
  NAND2XLTH U8 ( .A(A[2]), .B(B[2]), .Y(n4) );
  NAND2XLTH U9 ( .A(A[2]), .B(carry[2]), .Y(n3) );
  XOR2X1TH U10 ( .A(n2), .B(A[2]), .Y(SUM[2]) );
endmodule


module add_33_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_33_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7;
  wire   [5:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX4TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1TH U2 ( .A(A[6]), .B(B[6]), .Y(n6) );
  CLKXOR2X1TH U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2XLTH U4 ( .A(B[5]), .B(A[5]), .Y(n2) );
  XOR2X1TH U5 ( .A(n2), .B(carry[5]), .Y(SUM[5]) );
  NAND2XLTH U6 ( .A(carry[5]), .B(B[5]), .Y(n4) );
  NAND2XLTH U7 ( .A(carry[5]), .B(A[5]), .Y(n3) );
  NAND2XLTH U8 ( .A(A[5]), .B(B[5]), .Y(n5) );
  AND3X2 U9 ( .A(n3), .B(n4), .C(n5), .Y(n7) );
  XNOR2X4 U10 ( .A(n7), .B(n6), .Y(SUM[6]) );
endmodule


module add_33_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_33_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n7, n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXLTH U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(n7) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  NAND2X2TH U1 ( .A(n4), .B(n5), .Y(SUM[0]) );
  NAND2XLTH U2 ( .A(B[0]), .B(n3), .Y(n4) );
  NAND2XLTH U3 ( .A(n2), .B(A[0]), .Y(n5) );
  INVXLTH U4 ( .A(B[0]), .Y(n2) );
  INVXLTH U5 ( .A(A[0]), .Y(n3) );
  AND2XLTH U6 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKBUFX40 U7 ( .A(n7), .Y(SUM[1]) );
endmodule


module add_33_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  NAND2X4 U1 ( .A(n4), .B(n5), .Y(SUM[0]) );
  NAND2XL U2 ( .A(B[0]), .B(n3), .Y(n4) );
  NAND2X5 U3 ( .A(n2), .B(A[0]), .Y(n5) );
  INVX2TH U4 ( .A(B[0]), .Y(n2) );
  INVXLTH U5 ( .A(A[0]), .Y(n3) );
  AND2XLTH U6 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_33 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n21, n22, n23;

  add_33_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n23, 
        temp1_1_, temp1_0_}), .B(in2), .SUM(out3) );
  add_33_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_33_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n23, 
        temp1_1_, temp1_0_}), .B({in3[6], n22, in3[4:3], n21, in3[1:0]}), 
        .SUM(out2) );
  add_33_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n23, 
        temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_33_DW01_add_4 add_30 ( .A(in2), .B({in3[6], n22, in3[4:3], n21, in3[1:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_33_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX1TH U1 ( .A(in3[2]), .Y(n21) );
  CLKBUFX40 U2 ( .A(in3[5]), .Y(n22) );
  CLKBUFX40 U3 ( .A(temp1_2_), .Y(n23) );
endmodule


module tc_sm_135 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n28) );
  XNOR2XLTH U7 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(n31), .Y(n24) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(n31), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXLTH U11 ( .A(in[5]), .Y(n25) );
  INVXLTH U12 ( .A(in[4]), .Y(n26) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n27) );
  CLKBUFX1TH U14 ( .A(n31), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U16 ( .A0(n24), .A1(n12), .B0(n31), .B1(n29), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U17 ( .A0(n24), .A1(n10), .B0(n31), .B1(n28), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U18 ( .A0(n9), .A1(n27), .B0(n31), .Y(n7) );
  OAI211XLTH U19 ( .A0(n31), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n27), .A1N(n9), .B0(n31), .Y(n13) );
  CLKBUFX40 U21 ( .A(in[6]), .Y(n31) );
endmodule


module tc_sm_134 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n20, n21, n22, n23, n24, n25,
         n26;

  OAI33X2 U3 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n22), .B2(n23), .Y(n8) );
  OAI21X1 U4 ( .A0(in[3]), .A1(n20), .B0(in[6]), .Y(n13) );
  OAI211XLTH U5 ( .A0(in[6]), .A1(n24), .B0(n7), .C0(n18), .Y(out[3]) );
  BUFX10 U6 ( .A(n8), .Y(n18) );
  OAI221XL U7 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n25), .C0(n18), .Y(out[2])
         );
  OAI221XL U8 ( .A0(n21), .A1(n12), .B0(in[6]), .B1(n26), .C0(n18), .Y(out[1])
         );
  INVX2TH U9 ( .A(in[4]), .Y(n23) );
  INVXLTH U10 ( .A(in[6]), .Y(n21) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U12 ( .A(n9), .Y(n20) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U14 ( .A(n25), .B(n11), .Y(n10) );
  OAI21XLTH U15 ( .A0(n9), .A1(n24), .B0(in[6]), .Y(n7) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  INVX2 U17 ( .A(in[5]), .Y(n22) );
  INVXLTH U18 ( .A(in[3]), .Y(n24) );
  NOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U20 ( .A(in[2]), .Y(n25) );
  INVXLTH U21 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U22 ( .A(in[0]), .B(in[1]), .Y(n12) );
endmodule


module tc_sm_133 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n20, n21, n22, n23, n24, n25,
         n27;

  BUFX8 U3 ( .A(n8), .Y(n18) );
  OAI2BB1X2 U4 ( .A0N(n23), .A1N(n9), .B0(n27), .Y(n13) );
  OAI221XL U5 ( .A0(n20), .A1(n12), .B0(n27), .B1(n25), .C0(n18), .Y(out[1])
         );
  OAI221XL U6 ( .A0(n20), .A1(n10), .B0(n27), .B1(n24), .C0(n18), .Y(out[2])
         );
  OAI211XL U7 ( .A0(n27), .A1(n23), .B0(n7), .C0(n18), .Y(out[3]) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U10 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n12) );
  CLKBUFX1TH U12 ( .A(n27), .Y(out[4]) );
  XNOR2XLTH U13 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U15 ( .A(in[2]), .Y(n24) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  INVX4 U17 ( .A(in[5]), .Y(n21) );
  INVXLTH U18 ( .A(n27), .Y(n20) );
  OAI21XLTH U19 ( .A0(n9), .A1(n23), .B0(n27), .Y(n7) );
  OAI33X4 U20 ( .A0(in[4]), .A1(n27), .A2(in[5]), .B0(n13), .B1(n21), .B2(n22), 
        .Y(n8) );
  INVXL U21 ( .A(in[4]), .Y(n22) );
  CLKBUFX40 U22 ( .A(in[6]), .Y(n27) );
endmodule


module tc_sm_132 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n19, n20, n21, n23, n24, n25,
         n26, n27, n28;

  INVX2TH U3 ( .A(in[5]), .Y(n25) );
  BUFX10 U4 ( .A(n8), .Y(n18) );
  OR3XLTH U5 ( .A(n19), .B(n20), .C(n21), .Y(out[1]) );
  OAI221X1TH U6 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n23), .C0(n18), .Y(
        out[2]) );
  NOR2XLTH U7 ( .A(n24), .B(n12), .Y(n19) );
  NOR2XLTH U8 ( .A(in[6]), .B(n28), .Y(n20) );
  INVXLTH U9 ( .A(n18), .Y(n21) );
  INVXL U10 ( .A(in[6]), .Y(n24) );
  XNOR2X1TH U11 ( .A(in[0]), .B(in[1]), .Y(n12) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n27) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVX2TH U14 ( .A(in[4]), .Y(n26) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U16 ( .A(in[1]), .Y(n28) );
  XNOR2XLTH U17 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n18), .Y(out[3]) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  OAI21XLTH U21 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  OAI2BB1X4 U22 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
  INVXLTH U23 ( .A(in[2]), .Y(n23) );
  OAI33X4 U24 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
endmodule


module total_3_test_14 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n4, n5, n40, n41, n42, n49, n50, n51, n52, n53, n54, n55, n56;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_135 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_134 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_133 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_132 sm_tc_4 ( .out(in1), .in(in) );
  add_33 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_135 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_134 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_133 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_132 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up3[3]) );
  SDFFRQX1TH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n52), .CK(clk), .RN(n4), .Q(
        up1[0]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up2[3]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n53), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRQX1TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n53), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRQX2TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n53), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n56), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n56), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  SDFFRQX4TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n55), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n5) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n4) );
  SDFFRX4 h_reg ( .D(w5_4_), .SI(test_si), .SE(n52), .CK(clk), .RN(n5), .Q(h)
         );
  SDFFRHQX8 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n53), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up1[1]) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n55), .CK(clk), .RN(n4), 
        .Q(up1[2]) );
  INVXLTH U37 ( .A(test_se), .Y(n40) );
  INVXLTH U38 ( .A(n40), .Y(n41) );
  INVXLTH U39 ( .A(n40), .Y(n42) );
  DLY1X1TH U40 ( .A(n54), .Y(n49) );
  INVXLTH U41 ( .A(n49), .Y(n50) );
  INVXLTH U42 ( .A(n49), .Y(n51) );
  DLY1X1TH U43 ( .A(n41), .Y(n52) );
  DLY1X1TH U44 ( .A(n42), .Y(n53) );
  INVXLTH U45 ( .A(n41), .Y(n54) );
  INVXLTH U46 ( .A(n49), .Y(n55) );
  INVXLTH U47 ( .A(n49), .Y(n56) );
endmodule


module sm_tc_131 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n21, n22, n25, n26;

  XNOR2X2 U2 ( .A(n7), .B(n25), .Y(n4) );
  CLKBUFX2TH U3 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X4 U4 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  INVX4 U5 ( .A(n17), .Y(n22) );
  OAI2BB2XLTH U6 ( .B0(n22), .B1(n4), .A0N(n25), .A1N(n22), .Y(out[3]) );
  XNOR2X1TH U7 ( .A(n21), .B(n8), .Y(n5) );
  OAI22XL U8 ( .A0(n17), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  AOI31X1 U9 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  INVX2TH U10 ( .A(in[2]), .Y(n21) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  NOR2X6 U12 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[5]) );
  BUFX2 U14 ( .A(in[4]), .Y(n17) );
  NAND2XLTH U15 ( .A(n8), .B(n21), .Y(n7) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX40 U16 ( .A(in[3]), .Y(n25) );
  AOI21X8 U18 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n26) );
  CLKINVX40 U19 ( .A(n26), .Y(n6) );
endmodule


module sm_tc_130 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n19, n23, n26;

  OAI2BB2X2TH U2 ( .B0(n19), .B1(n6), .A0N(in[1]), .A1N(n19), .Y(out[1]) );
  NOR2X4 U3 ( .A(in[1]), .B(n26), .Y(n8) );
  INVX2TH U4 ( .A(in[4]), .Y(n19) );
  AO21XLTH U5 ( .A0(n26), .A1(in[1]), .B0(n8), .Y(n6) );
  XNOR2X1TH U6 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI22XL U7 ( .A0(in[4]), .A1(n23), .B0(n19), .B1(n5), .Y(out[2]) );
  CLKBUFX2TH U9 ( .A(n26), .Y(out[0]) );
  INVX2 U10 ( .A(in[2]), .Y(n23) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  NAND2XLTH U12 ( .A(n8), .B(n23), .Y(n7) );
  NOR2BXLTH U13 ( .AN(n6), .B(n26), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2X1TH U15 ( .B0(n19), .B1(n4), .A0N(in[3]), .A1N(n19), .Y(out[3]) );
  AOI31X2TH U16 ( .A0(n3), .A1(n4), .A2(n5), .B0(n19), .Y(out[4]) );
  CLKBUFX40 U8 ( .A(in[0]), .Y(n26) );
  XOR2X1 U17 ( .A(in[2]), .B(n8), .Y(n5) );
endmodule


module sm_tc_129 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n6, n8, n25, n26, n27, n31, n32, n35, n36, n37, n38;

  NOR2X4 U2 ( .A(n37), .B(in[0]), .Y(n8) );
  OR2X2 U3 ( .A(n31), .B(n38), .Y(n27) );
  INVX4 U4 ( .A(n25), .Y(n31) );
  OAI2BB2X1 U5 ( .B0(n31), .B1(n4), .A0N(in[3]), .A1N(n31), .Y(out[3]) );
  AOI31X2 U6 ( .A0(n3), .A1(n4), .A2(n38), .B0(n31), .Y(out[4]) );
  OAI2BB2X2 U7 ( .B0(n31), .B1(n6), .A0N(n37), .A1N(n31), .Y(out[1]) );
  CLKBUFX1TH U9 ( .A(in[4]), .Y(n25) );
  INVX1TH U11 ( .A(in[2]), .Y(n32) );
  OR2XLTH U12 ( .A(n25), .B(n35), .Y(n26) );
  CLKNAND2X2TH U13 ( .A(n26), .B(n27), .Y(out[2]) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U16 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[6]) );
  NOR2BXLTH U18 ( .AN(n6), .B(in[0]), .Y(n3) );
  AO21XLTH U19 ( .A0(in[0]), .A1(n37), .B0(n8), .Y(n6) );
  CLKBUFX40 U8 ( .A(n32), .Y(n35) );
  XNOR2X1 U10 ( .A(n35), .B(n8), .Y(n38) );
  XOR2X1 U15 ( .A(n36), .B(in[3]), .Y(n4) );
  CLKAND2X12 U20 ( .A(n35), .B(n8), .Y(n36) );
  CLKBUFX40 U21 ( .A(in[1]), .Y(n37) );
endmodule


module sm_tc_128 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  AOI31X2 U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  CLKBUFX1TH U3 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1TH U4 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U5 ( .A(n8), .B(n21), .Y(n7) );
  OAI2BB2X1TH U6 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  CLKINVX1TH U7 ( .A(n18), .Y(out[5]) );
  NOR2X6TH U8 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX2TH U9 ( .A(in[4]), .Y(n22) );
  OAI2BB2X2TH U10 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n21) );
  INVXLTH U12 ( .A(out[4]), .Y(n18) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI22X1TH U14 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  INVXLTH U15 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U16 ( .A(n21), .B(n8), .Y(n5) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_32_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR3X2 U3 ( .A(A[6]), .B(n3), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
  CLKINVX40 U5 ( .A(B[6]), .Y(n3) );
endmodule


module add_32_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [6:2] carry;

  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X12 U1 ( .A(n6), .B(carry[6]), .Y(SUM[6]) );
  XOR2X1 U2 ( .A(n2), .B(carry[5]), .Y(SUM[5]) );
  XOR2X1 U3 ( .A(B[5]), .B(A[5]), .Y(n2) );
  NAND2XLTH U4 ( .A(A[5]), .B(B[5]), .Y(n5) );
  NAND2XLTH U5 ( .A(carry[5]), .B(B[5]), .Y(n4) );
  NAND3X2 U6 ( .A(n3), .B(n4), .C(n5), .Y(carry[6]) );
  AND2XLTH U7 ( .A(n8), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U8 ( .A(n8), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U9 ( .A(B[6]), .B(A[6]), .Y(n6) );
  NAND2XLTH U10 ( .A(carry[5]), .B(A[5]), .Y(n3) );
  INVXLTH U11 ( .A(B[0]), .Y(n7) );
  INVXLTH U12 ( .A(n7), .Y(n8) );
endmodule


module add_32_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_32_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n3;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR2X4TH U2 ( .A(n3), .B(carry[6]), .Y(SUM[6]) );
  XNOR2XLTH U3 ( .A(A[6]), .B(B[6]), .Y(n3) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_32_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(n2), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKINVX40 U4 ( .A(A[6]), .Y(n2) );
endmodule


module add_32_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2TH U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U2 ( .A(B[0]), .B(n3), .Y(n1) );
  DLY1X1TH U1 ( .A(n4), .Y(n2) );
  INVXLTH U3 ( .A(n5), .Y(n3) );
  XOR2X1 U4 ( .A(B[0]), .B(n5), .Y(n4) );
  CLKINVX40 U5 ( .A(n2), .Y(SUM[0]) );
  CLKINVX40 U6 ( .A(A[0]), .Y(n5) );
endmodule


module add_32 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;

  add_32_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n28, temp1_2_, 
        n23, temp1_0_}), .B({n26, in2[5:3], n18, n21, in2[0]}), .SUM(out3) );
  add_32_DW01_add_1 add_33 ( .A({temp2_6_, n22, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_32_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n28, temp1_2_, 
        n23, temp1_0_}), .B({in3[6:2], n24, n27}), .SUM(out2) );
  add_32_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n28, temp1_2_, 
        n23, temp1_0_}), .B({temp2_6_, n22, temp2_4_, temp2_3_, temp2_2_, n19, 
        temp2_0_}), .SUM(out) );
  add_32_DW01_add_4 add_30 ( .A({n25, in2[5:3], n18, n21, in2[0]}), .B({
        in3[6:2], n24, n27}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}) );
  add_32_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  INVX2TH U1 ( .A(n20), .Y(n21) );
  INVX2 U2 ( .A(in2[1]), .Y(n20) );
  BUFX2TH U3 ( .A(in2[2]), .Y(n18) );
  CLKBUFX1TH U4 ( .A(temp2_1_), .Y(n19) );
  CLKBUFX40 U5 ( .A(temp2_5_), .Y(n22) );
  CLKBUFX40 U6 ( .A(temp1_1_), .Y(n23) );
  CLKBUFX40 U13 ( .A(in3[1]), .Y(n24) );
  DLY1X1TH U14 ( .A(in2[6]), .Y(n25) );
  DLY1X1TH U15 ( .A(in2[6]), .Y(n26) );
  CLKBUFX40 U16 ( .A(in3[0]), .Y(n27) );
  CLKBUFX40 U17 ( .A(temp1_3_), .Y(n28) );
endmodule


module tc_sm_131 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31, n33;

  BUFX2 U3 ( .A(n33), .Y(out[4]) );
  NOR3X1TH U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U5 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U6 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U7 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U8 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(n33), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n28) );
  INVXLTH U12 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n29) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(n33), .Y(n26) );
  OAI21XLTH U16 ( .A0(n9), .A1(n29), .B0(n33), .Y(n7) );
  OAI221XLTH U17 ( .A0(n26), .A1(n12), .B0(n33), .B1(n31), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U18 ( .A0(n26), .A1(n10), .B0(n33), .B1(n30), .C0(n8), .Y(out[2])
         );
  OAI211XLTH U19 ( .A0(n33), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(n33), .Y(n13) );
  CLKBUFX40 U21 ( .A(in[6]), .Y(n33) );
endmodule


module tc_sm_130 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n20, n21, n22, n23, n25, n26;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(n26), .Y(n11) );
  OAI211XL U3 ( .A0(in[6]), .A1(n21), .B0(n5), .C0(n6), .Y(out[3]) );
  AOI21X8 U4 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n6) );
  INVXLTH U5 ( .A(in[6]), .Y(n20) );
  OAI221X1 U6 ( .A0(n25), .A1(n10), .B0(in[6]), .B1(n23), .C0(n6), .Y(out[1])
         );
  OAI221X2TH U8 ( .A0(n20), .A1(n8), .B0(in[6]), .B1(n22), .C0(n6), .Y(out[2])
         );
  AOI2BB1X2TH U9 ( .A0N(n26), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U11 ( .A(in[6]), .Y(out[4]) );
  XOR2XLTH U12 ( .A(in[0]), .B(n23), .Y(n10) );
  INVXLTH U13 ( .A(in[1]), .Y(n23) );
  INVXLTH U14 ( .A(in[2]), .Y(n22) );
  XOR2XLTH U15 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n9) );
  INVXLTH U17 ( .A(in[3]), .Y(n21) );
  OAI21XLTH U18 ( .A0(n7), .A1(n21), .B0(in[6]), .Y(n5) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  INVXLTH U20 ( .A(in[6]), .Y(n25) );
  CLKBUFX40 U21 ( .A(in[5]), .Y(n26) );
endmodule


module tc_sm_129 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n20, n21, n22, n24, n25, n26, n27,
         n28, n29, n31;

  BUFX6 U3 ( .A(n8), .Y(n20) );
  OAI211XLTH U5 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n20), .Y(out[3]) );
  OR2XLTH U6 ( .A(n24), .B(n12), .Y(n21) );
  OR2XLTH U7 ( .A(in[6]), .B(n29), .Y(n22) );
  NAND2BXL U8 ( .AN(in[0]), .B(n20), .Y(out[0]) );
  OAI221XL U9 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n20), .Y(out[2])
         );
  OAI2BB1X4 U10 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
  INVXLTH U11 ( .A(in[6]), .Y(n24) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n27) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U14 ( .A(n28), .B(n11), .Y(n10) );
  INVXLTH U15 ( .A(in[2]), .Y(n28) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI21XLTH U17 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U18 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U19 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVX2 U21 ( .A(in[5]), .Y(n25) );
  OAI33X4 U22 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXL U23 ( .A(in[4]), .Y(n26) );
  AND3X8 U4 ( .A(n21), .B(n22), .C(n20), .Y(n31) );
  CLKINVX40 U24 ( .A(n31), .Y(out[1]) );
endmodule


module tc_sm_128 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n21, n23, n24, n25, n26;

  AOI21BX4TH U3 ( .A0(in[6]), .A1(n11), .B0N(n21), .Y(n6) );
  OAI21BX4TH U4 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n21) );
  OAI2B11X2TH U5 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  INVXLTH U6 ( .A(in[6]), .Y(n23) );
  NOR3X1TH U7 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  INVXLTH U8 ( .A(in[2]), .Y(n25) );
  XOR2XLTH U9 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U10 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI211XLTH U11 ( .A0(in[6]), .A1(n24), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI21XLTH U12 ( .A0(n7), .A1(n24), .B0(in[6]), .Y(n5) );
  INVXLTH U13 ( .A(in[3]), .Y(n24) );
  XOR2XLTH U14 ( .A(in[0]), .B(n26), .Y(n10) );
  INVXLTH U15 ( .A(in[1]), .Y(n26) );
  CLKBUFX1TH U16 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  OAI221XLTH U18 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n26), .C0(n6), .Y(
        out[1]) );
  OAI221XLTH U19 ( .A0(n23), .A1(n8), .B0(in[6]), .B1(n25), .C0(n6), .Y(out[2]) );
endmodule


module total_3_test_15 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n63, n64, w5_4_, n4, n5, n40, n48, n49, n50, n51, n52, n53, n54, n55;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_131 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_130 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_129 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_128 sm_tc_4 ( .out(in1), .in(in) );
  add_32 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_131 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_130 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_129 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_128 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXL up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(n64) );
  SDFFRQXL up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(n63) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n49), .CK(clk), .RN(n5), .Q(
        up1[0]) );
  SDFFRQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n54), .CK(clk), .RN(n4), 
        .Q(up1[4]) );
  SDFFRQX2 up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n55), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n55), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRQX1TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up2[4]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n5) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n4) );
  SDFFRX4 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n54), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up1[1]) );
  SDFFRX4 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  SDFFRX4 h_reg ( .D(w5_4_), .SI(test_si), .SE(n49), .CK(clk), .RN(n5), .Q(h)
         );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  INVXLTH U37 ( .A(n53), .Y(n40) );
  DLY1X1TH U38 ( .A(n63), .Y(up1[2]) );
  DLY1X1TH U39 ( .A(n53), .Y(n48) );
  INVXLTH U40 ( .A(n48), .Y(n49) );
  INVXLTH U41 ( .A(n48), .Y(n50) );
  DLY1X1TH U42 ( .A(n40), .Y(n51) );
  DLY1X1TH U43 ( .A(test_se), .Y(n52) );
  INVXLTH U44 ( .A(test_se), .Y(n53) );
  INVXLTH U45 ( .A(n48), .Y(n54) );
  INVXLTH U46 ( .A(n48), .Y(n55) );
  DLY1X1TH U47 ( .A(n64), .Y(up3[3]) );
endmodule


module sm_tc_127 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n20, n21, n24, n25, n26;

  OAI2BB2X1 U2 ( .B0(n21), .B1(n4), .A0N(in[3]), .A1N(n21), .Y(out[3]) );
  INVX6 U5 ( .A(in[4]), .Y(n21) );
  AOI31X1 U6 ( .A0(n3), .A1(n4), .A2(n5), .B0(n21), .Y(out[4]) );
  OAI22XL U7 ( .A0(in[4]), .A1(n20), .B0(n21), .B1(n5), .Y(out[2]) );
  XNOR2X1 U8 ( .A(n20), .B(n8), .Y(n5) );
  AO21X1 U10 ( .A0(n25), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X6 U11 ( .A(in[1]), .B(n25), .Y(n8) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[6]) );
  INVX1TH U13 ( .A(in[2]), .Y(n20) );
  NOR2BXLTH U14 ( .AN(n6), .B(n25), .Y(n3) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  BUFX2TH U16 ( .A(n25), .Y(out[0]) );
  XOR2X1 U3 ( .A(n24), .B(in[3]), .Y(n4) );
  CLKAND2X12 U4 ( .A(n8), .B(n20), .Y(n24) );
  CLKBUFX40 U9 ( .A(in[0]), .Y(n25) );
  AO2B2X4 U17 ( .B0(in[1]), .B1(n21), .A0(n26), .A1N(n6), .Y(out[1]) );
  CLKINVX40 U18 ( .A(n21), .Y(n26) );
endmodule


module sm_tc_126 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n30, n31, n33, n34, n35, n40, n41, n44, n45;

  AO21X1 U2 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  BUFX3 U3 ( .A(in[0]), .Y(out[0]) );
  NOR2X6 U4 ( .A(in[1]), .B(in[0]), .Y(n8) );
  BUFX10 U5 ( .A(in[4]), .Y(n30) );
  NAND2X2 U9 ( .A(n34), .B(n35), .Y(n4) );
  AND3XL U10 ( .A(n3), .B(n4), .C(n5), .Y(n31) );
  INVX2 U11 ( .A(n30), .Y(n40) );
  OAI2BB2X2TH U13 ( .B0(n40), .B1(n4), .A0N(in[3]), .A1N(n40), .Y(out[3]) );
  INVX1TH U14 ( .A(in[2]), .Y(n41) );
  CLKNAND2X2TH U15 ( .A(n7), .B(in[3]), .Y(n34) );
  CLKNAND2X4 U17 ( .A(n44), .B(n33), .Y(n35) );
  XNOR2X1TH U18 ( .A(n41), .B(n8), .Y(n5) );
  INVXLTH U19 ( .A(in[3]), .Y(n33) );
  INVXLTH U20 ( .A(n45), .Y(out[6]) );
  INVXLTH U21 ( .A(n45), .Y(out[5]) );
  NOR2BXLTH U22 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2B2X2 U6 ( .A1N(in[1]), .A0(n30), .B0(n40), .B1(n6), .Y(out[1]) );
  AND2X8 U7 ( .A(n8), .B(n41), .Y(n44) );
  CLKINVX40 U8 ( .A(n44), .Y(n7) );
  OAI2B2X2 U12 ( .A1N(n30), .A0(n5), .B0(n30), .B1(n41), .Y(out[2]) );
  NAND2BX8 U16 ( .AN(n31), .B(n30), .Y(n45) );
  CLKINVX40 U23 ( .A(n45), .Y(out[4]) );
endmodule


module sm_tc_125 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n23, n24, n28, n29;

  BUFX2 U2 ( .A(out[6]), .Y(out[4]) );
  CLKBUFX2TH U3 ( .A(out[6]), .Y(out[5]) );
  AOI31X2 U4 ( .A0(n3), .A1(n4), .A2(n5), .B0(n28), .Y(out[6]) );
  BUFX4 U5 ( .A(in[4]), .Y(n24) );
  AO21X2 U6 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2X4 U7 ( .B0(n28), .B1(n6), .A0N(in[1]), .A1N(n28), .Y(out[1]) );
  NOR2X6 U8 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X1TH U9 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U10 ( .A(n8), .B(n29), .Y(n7) );
  NOR2XLTH U11 ( .A(n24), .B(n29), .Y(n22) );
  NOR2X1 U12 ( .A(n28), .B(n5), .Y(n23) );
  OR2X2 U13 ( .A(n22), .B(n23), .Y(out[2]) );
  INVX4 U14 ( .A(n24), .Y(n28) );
  OAI2BB2X1 U15 ( .B0(n28), .B1(n4), .A0N(in[3]), .A1N(n28), .Y(out[3]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX2 U17 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1TH U18 ( .A(n29), .B(n8), .Y(n5) );
  INVX2 U19 ( .A(in[2]), .Y(n29) );
endmodule


module sm_tc_124 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  CLKBUFX1TH U2 ( .A(in[0]), .Y(out[0]) );
  NOR2X3TH U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI22X1TH U4 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  OAI2BB2X2TH U5 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  INVXLTH U6 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U7 ( .A(n7), .B(in[3]), .Y(n4) );
  XNOR2X1TH U8 ( .A(n21), .B(n8), .Y(n5) );
  CLKINVX1TH U9 ( .A(in[2]), .Y(n21) );
  CLKINVX2TH U10 ( .A(in[4]), .Y(n22) );
  OAI2BB2X1TH U11 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  AOI31X2TH U12 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U14 ( .A(out[4]), .Y(n18) );
  INVXLTH U15 ( .A(n18), .Y(out[5]) );
  NAND2XLTH U16 ( .A(n8), .B(n21), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_31_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_31_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_31_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_31_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_31_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_31_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_31 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n16, n17, n18;

  add_31_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n18, temp1_0_}), .B(in2), .SUM(out3) );
  add_31_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, n16}), .B(in), .SUM(out1) );
  add_31_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n18, temp1_0_}), .B(in3), .SUM(out2) );
  add_31_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n18, n17}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, n16}), .SUM(out) );
  add_31_DW01_add_4 add_30 ( .A(in2), .B(in3), .SUM({temp2_6_, temp2_5_, 
        temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_31_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2 U1 ( .A(temp2_0_), .Y(n16) );
  CLKBUFX1TH U2 ( .A(temp1_0_), .Y(n17) );
  CLKBUFX40 U3 ( .A(temp1_1_), .Y(n18) );
endmodule


module tc_sm_127 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n28) );
  XNOR2XLTH U7 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(in[6]), .Y(n24) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n26) );
  INVXLTH U12 ( .A(in[5]), .Y(n25) );
  OAI21XLTH U13 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  CLKINVX1TH U14 ( .A(in[3]), .Y(n27) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  OAI221XLTH U16 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(
        out[2]) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_126 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n23, n24, n25, n27, n28, n29,
         n30, n31, n32;

  OAI211XL U4 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221XL U6 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[1])
         );
  OAI221X2TH U7 ( .A0(n29), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[2]) );
  NAND2BXLTH U8 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n23) );
  INVXLTH U10 ( .A(in[6]), .Y(n20) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U12 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U14 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U16 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  INVX2 U18 ( .A(in[5]), .Y(n21) );
  INVXLTH U19 ( .A(in[2]), .Y(n24) );
  AOI33X4 U3 ( .A0(n28), .A1(n29), .A2(n21), .B0(n32), .B1(n30), .B2(n31), .Y(
        n27) );
  CLKINVX40 U5 ( .A(n27), .Y(n8) );
  CLKINVX40 U20 ( .A(in[4]), .Y(n28) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n29) );
  CLKINVX40 U22 ( .A(n21), .Y(n30) );
  CLKINVX40 U23 ( .A(n28), .Y(n31) );
  AOI21BX4 U24 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n32) );
endmodule


module tc_sm_125 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n35, n37, n38, n39, n40;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[5]), .C0(in[4]), .Y(n11) );
  OAI221XL U3 ( .A0(n37), .A1(n10), .B0(in[6]), .B1(n40), .C0(n6), .Y(out[1])
         );
  INVXL U4 ( .A(in[6]), .Y(n37) );
  AOI21BX4 U5 ( .A0(in[6]), .A1(n11), .B0N(n35), .Y(n6) );
  OAI21XLTH U6 ( .A0(n7), .A1(n38), .B0(in[6]), .Y(n5) );
  INVXLTH U8 ( .A(in[3]), .Y(n38) );
  NAND2BXLTH U9 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  INVXLTH U10 ( .A(in[2]), .Y(n39) );
  XOR2XLTH U11 ( .A(in[2]), .B(n9), .Y(n8) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U13 ( .A(in[1]), .Y(n40) );
  OAI21BX1 U14 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n35) );
  NOR3X1TH U15 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  OAI221XLTH U16 ( .A0(n37), .A1(n8), .B0(in[6]), .B1(n39), .C0(n6), .Y(out[2]) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n9) );
  XOR2XLTH U18 ( .A(in[0]), .B(n40), .Y(n10) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n38), .B0(n5), .C0(n6), .Y(out[3]) );
endmodule


module tc_sm_124 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n11, n12, n13, n36, n37, n38, n39, n41, n42, n43;

  NOR3X4 U3 ( .A(in[5]), .B(in[6]), .C(in[4]), .Y(n5) );
  OAI221XL U4 ( .A0(n36), .A1(n12), .B0(in[6]), .B1(n39), .C0(n41), .Y(out[1])
         );
  AOI21X1 U5 ( .A0(n5), .A1(n37), .B0(n6), .Y(out[3]) );
  AOI31X2 U7 ( .A0(in[5]), .A1(n13), .A2(in[4]), .B0(n36), .Y(n8) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n37) );
  NAND2XLTH U9 ( .A(n37), .B(n7), .Y(n13) );
  CLKINVX3TH U10 ( .A(in[6]), .Y(n36) );
  NOR3X4TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  XOR2XLTH U14 ( .A(in[0]), .B(n39), .Y(n12) );
  INVXLTH U15 ( .A(in[1]), .Y(n39) );
  OAI21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(in[2]), .Y(n11) );
  AOI32XLTH U18 ( .A0(in[6]), .A1(n38), .A2(n11), .B0(in[2]), .B1(n36), .Y(n9)
         );
  INVXLTH U19 ( .A(n7), .Y(n38) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n41), .Y(out[0]) );
  AOI2BB1X4 U6 ( .A0N(in[6]), .A1N(n5), .B0(n8), .Y(n41) );
  AND2X8 U11 ( .A(n9), .B(n41), .Y(n42) );
  CLKINVX40 U16 ( .A(n42), .Y(out[2]) );
  NOR4BBX4 U21 ( .AN(n43), .BN(in[6]), .C(n8), .D(n37), .Y(n6) );
  CLKINVX40 U22 ( .A(n7), .Y(n43) );
endmodule


module total_3_test_16 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n4, n5, n6, n7, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_127 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_126 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_125 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_124 sm_tc_4 ( .out(in1), .in(in) );
  add_31 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2({b1[6:2], n54, b1[0]}), .in3({c1[6:1], n5}), .in(in1) );
  tc_sm_127 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_126 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_125 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_124 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n49), .CK(clk), .RN(n7), .Q(
        h) );
  SDFFRQXLTH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up2[1]) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n47), .CK(clk), .RN(n6), 
        .Q(up1[4]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n52), .CK(clk), .RN(n6), 
        .Q(up2[2]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up3[2]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up2[3]) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n45), .CK(clk), .RN(n6), 
        .Q(up3[3]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n53), .CK(clk), .RN(n6), 
        .Q(up2[0]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up3[0]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n45), .CK(clk), .RN(n7), 
        .Q(up1[3]) );
  SDFFRQX1TH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n53), .CK(clk), .RN(n6), 
        .Q(up1[1]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up3[4]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n47), .CK(clk), .RN(n7), 
        .Q(up1[2]) );
  SDFFRQX2 up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n52), .CK(clk), .RN(n6), .Q(
        up1[0]) );
  INVX6 U3 ( .A(c1[0]), .Y(n4) );
  CLKINVX16 U4 ( .A(n4), .Y(n5) );
  CLKBUFX4TH U5 ( .A(rst), .Y(n6) );
  CLKBUFX1TH U6 ( .A(rst), .Y(n7) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up3[1]) );
  DLY1X1TH U39 ( .A(n46), .Y(n44) );
  INVXLTH U40 ( .A(n46), .Y(n45) );
  DLY1X1TH U41 ( .A(n50), .Y(n46) );
  INVXLTH U42 ( .A(n46), .Y(n47) );
  INVXLTH U43 ( .A(n50), .Y(n48) );
  DLY1X1TH U44 ( .A(test_se), .Y(n49) );
  INVXLTH U45 ( .A(test_se), .Y(n50) );
  INVXLTH U46 ( .A(n44), .Y(n51) );
  INVXLTH U47 ( .A(n44), .Y(n52) );
  INVXLTH U48 ( .A(n46), .Y(n53) );
  CLKBUFX40 U49 ( .A(b1[1]), .Y(n54) );
endmodule


module sm_tc_123 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n18, n22, n23, n25, n26, n27, n28;

  XNOR2X2 U2 ( .A(n23), .B(n8), .Y(n5) );
  CLKBUFX4 U3 ( .A(in[0]), .Y(out[0]) );
  INVX4 U6 ( .A(in[4]), .Y(n22) );
  AND2X2 U7 ( .A(n18), .B(in[4]), .Y(out[6]) );
  INVX2TH U8 ( .A(in[2]), .Y(n23) );
  CLKBUFX2 U9 ( .A(out[6]), .Y(out[4]) );
  AO21X2 U11 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NAND3XL U13 ( .A(n3), .B(n26), .C(n5), .Y(n18) );
  NOR2BXL U14 ( .AN(n6), .B(out[0]), .Y(n3) );
  OAI2BB2XL U15 ( .B0(n25), .B1(n4), .A0N(in[3]), .A1N(n25), .Y(out[3]) );
  OAI2BB2X4TH U16 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U17 ( .A(out[6]), .Y(out[5]) );
  INVX4 U4 ( .A(in[4]), .Y(n25) );
  XNOR2X1 U5 ( .A(n28), .B(in[3]), .Y(n26) );
  OR2X8 U10 ( .A(in[1]), .B(out[0]), .Y(n27) );
  CLKINVX40 U12 ( .A(n27), .Y(n8) );
  AO2B2BX4 U18 ( .A0(n25), .A1N(n23), .B0(in[4]), .B1N(n5), .Y(out[2]) );
  XNOR2X1 U19 ( .A(n28), .B(in[3]), .Y(n4) );
  CLKNAND2X12 U20 ( .A(n8), .B(n23), .Y(n28) );
endmodule


module sm_tc_122 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n30, n31, n33, n36, n37;

  INVX2 U2 ( .A(in[2]), .Y(n36) );
  AOI31X2 U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n37), .Y(out[4]) );
  XNOR2X4 U4 ( .A(n36), .B(n8), .Y(n5) );
  BUFX2 U5 ( .A(in[4]), .Y(n30) );
  CLKBUFX2TH U6 ( .A(in[1]), .Y(n31) );
  OAI22X1TH U7 ( .A0(n30), .A1(n36), .B0(n37), .B1(n5), .Y(out[2]) );
  BUFX2 U8 ( .A(in[0]), .Y(out[0]) );
  AO21X1 U9 ( .A0(in[0]), .A1(n31), .B0(n8), .Y(n6) );
  CLKNAND2X2 U10 ( .A(n8), .B(n36), .Y(n7) );
  NOR2X4 U11 ( .A(n31), .B(in[0]), .Y(n8) );
  OAI2BB2X4TH U13 ( .B0(n37), .B1(n4), .A0N(in[3]), .A1N(n37), .Y(out[3]) );
  INVX2TH U14 ( .A(n30), .Y(n37) );
  XNOR2X2TH U15 ( .A(n7), .B(in[3]), .Y(n4) );
  INVXLTH U16 ( .A(out[4]), .Y(n33) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX1TH U18 ( .A(n33), .Y(out[5]) );
  INVXLTH U19 ( .A(n33), .Y(out[6]) );
  OAI2B2X2 U12 ( .A1N(n31), .A0(n30), .B0(n37), .B1(n6), .Y(out[1]) );
endmodule


module sm_tc_121 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n24, n25, n28, n29, n30;

  CLKNAND2X4 U2 ( .A(n28), .B(n24), .Y(n7) );
  BUFX5 U3 ( .A(in[0]), .Y(out[0]) );
  AO21X2 U4 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  XNOR2X2 U5 ( .A(n24), .B(n28), .Y(n5) );
  INVX4 U6 ( .A(in[4]), .Y(n25) );
  OAI2BB2X1 U7 ( .B0(n30), .B1(n4), .A0N(in[3]), .A1N(n30), .Y(out[3]) );
  XNOR2X4 U8 ( .A(n7), .B(in[3]), .Y(n4) );
  NOR2X4 U10 ( .A(in[1]), .B(out[0]), .Y(n8) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  OAI22X2TH U12 ( .A0(in[4]), .A1(n24), .B0(n30), .B1(n5), .Y(out[2]) );
  AOI31X2TH U13 ( .A0(n3), .A1(n4), .A2(n5), .B0(n30), .Y(out[4]) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  INVX2 U15 ( .A(in[2]), .Y(n24) );
  NOR2BXLTH U16 ( .AN(n6), .B(out[0]), .Y(n3) );
  AO2B2X4 U9 ( .B0(in[1]), .B1(n30), .A0(n29), .A1N(n6), .Y(out[1]) );
  CLKBUFX40 U17 ( .A(n8), .Y(n28) );
  CLKINVX40 U18 ( .A(n25), .Y(n29) );
  CLKINVX40 U19 ( .A(n29), .Y(n30) );
endmodule


module sm_tc_120 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n18, n19, n20, n24, n25;

  AOI31X2TH U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n25), .Y(out[6]) );
  NAND2XLTH U3 ( .A(n24), .B(n8), .Y(n19) );
  NAND2X2 U4 ( .A(n17), .B(n18), .Y(n20) );
  NAND2X2 U5 ( .A(n19), .B(n20), .Y(n5) );
  INVXL U6 ( .A(n24), .Y(n17) );
  INVXLTH U7 ( .A(n8), .Y(n18) );
  NOR2X4 U8 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI22X1 U9 ( .A0(in[4]), .A1(n24), .B0(n25), .B1(n5), .Y(out[2]) );
  CLKBUFX1TH U10 ( .A(in[0]), .Y(out[0]) );
  NAND2X1TH U11 ( .A(n8), .B(n24), .Y(n7) );
  OAI2BB2X2TH U12 ( .B0(n25), .B1(n4), .A0N(in[3]), .A1N(n25), .Y(out[3]) );
  CLKINVX2TH U13 ( .A(in[4]), .Y(n25) );
  CLKINVX1TH U14 ( .A(in[2]), .Y(n24) );
  OAI2BB2X2TH U15 ( .B0(n25), .B1(n6), .A0N(in[1]), .A1N(n25), .Y(out[1]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  XNOR2X1TH U17 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX1TH U18 ( .A(out[6]), .Y(out[4]) );
  CLKBUFX1TH U19 ( .A(out[6]), .Y(out[5]) );
  AO21XLTH U20 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_30_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR3X4TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_30_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_30_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_30_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_30_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [6:2] carry;

  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2TH U1_1 ( .A(B[1]), .B(n5), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  NAND2XL U1 ( .A(carry[3]), .B(B[3]), .Y(n2) );
  XOR2X1TH U2 ( .A(A[3]), .B(B[3]), .Y(n1) );
  NAND3X2 U3 ( .A(n2), .B(n3), .C(n4), .Y(carry[4]) );
  CLKXOR2X1TH U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U5 ( .A(B[0]), .B(A[0]), .Y(n5) );
  CLKXOR2X2TH U6 ( .A(n1), .B(carry[3]), .Y(SUM[3]) );
  NAND2XLTH U7 ( .A(B[3]), .B(A[3]), .Y(n4) );
  AND2X8 U8 ( .A(carry[3]), .B(A[3]), .Y(n6) );
  CLKINVX40 U9 ( .A(n6), .Y(n3) );
endmodule


module add_30_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2TH U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_30 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n27, n28, n29, n30;

  add_30_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, n29, temp1_3_, temp1_2_, 
        n28, temp1_0_}), .B(in2), .SUM(out3) );
  add_30_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_30_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, n29, temp1_3_, temp1_2_, 
        n28, temp1_0_}), .B({in3[6:4], n30, in3[2:0]}), .SUM(out2) );
  add_30_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, n29, temp1_3_, temp1_2_, 
        n28, temp1_0_}), .B({temp2_6_, temp2_5_, n27, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_30_DW01_add_4 add_30 ( .A(in2), .B({in3[6:4], n30, in3[2:0]}), .SUM({
        temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_})
         );
  add_30_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX1TH U1 ( .A(temp2_4_), .Y(n27) );
  CLKBUFX40 U2 ( .A(temp1_1_), .Y(n28) );
  CLKBUFX40 U3 ( .A(temp1_4_), .Y(n29) );
  CLKBUFX40 U4 ( .A(in3[3]), .Y(n30) );
endmodule


module tc_sm_123 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31, n33;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(n33), .A2(in[5]), .B0(n13), .B1(n27), .B2(n28), .Y(n8) );
  INVXLTH U10 ( .A(in[4]), .Y(n28) );
  INVXLTH U11 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(n33), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(n33), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(n33), .B1(n31), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(n33), .B1(n30), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(n33), .Y(n7) );
  OAI2BB1XLTH U19 ( .A0N(n29), .A1N(n9), .B0(n33), .Y(n13) );
  OAI211XLTH U20 ( .A0(n33), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  CLKBUFX40 U21 ( .A(in[6]), .Y(n33) );
endmodule


module tc_sm_122 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n6, n7, n8, n9, n10, n11, n19, n20, n22, n23, n24, n25, n26, n28, n29,
         n30, n31, n32;

  OAI221X2 U3 ( .A0(n28), .A1(n9), .B0(in[6]), .B1(n25), .C0(n7), .Y(out[2])
         );
  CLKINVX12 U4 ( .A(n19), .Y(n7) );
  CLKBUFX1TH U5 ( .A(in[6]), .Y(out[4]) );
  OAI221X1 U6 ( .A0(n28), .A1(n11), .B0(in[6]), .B1(n26), .C0(n7), .Y(out[1])
         );
  INVX1 U8 ( .A(in[6]), .Y(n22) );
  OA21X1 U9 ( .A0(n29), .A1(n8), .B0(in[6]), .Y(n20) );
  INVXLTH U10 ( .A(in[5]), .Y(n23) );
  NAND2XLTH U11 ( .A(n10), .B(n25), .Y(n8) );
  OAI2BB1XLTH U12 ( .A0N(n8), .A1N(in[3]), .B0(in[6]), .Y(n6) );
  NOR2XLTH U13 ( .A(in[1]), .B(n30), .Y(n10) );
  CLKINVX1TH U14 ( .A(in[2]), .Y(n25) );
  XNOR2XLTH U15 ( .A(n25), .B(n10), .Y(n9) );
  INVXLTH U16 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  AOI33X4 U18 ( .A0(n24), .A1(n28), .A2(n23), .B0(n20), .B1(in[5]), .B2(in[4]), 
        .Y(n19) );
  CLKINVX1 U19 ( .A(in[4]), .Y(n24) );
  CLKBUFX40 U7 ( .A(n22), .Y(n28) );
  INVXLTH U20 ( .A(n32), .Y(n29) );
  INVXLTH U21 ( .A(n31), .Y(n30) );
  NAND2X8 U22 ( .A(n31), .B(n7), .Y(out[0]) );
  CLKINVX40 U23 ( .A(in[0]), .Y(n31) );
  OAI211X4 U24 ( .A0(n32), .A1(in[6]), .B0(n6), .C0(n7), .Y(out[3]) );
  CLKINVX40 U25 ( .A(in[3]), .Y(n32) );
endmodule


module tc_sm_121 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n20, n21, n22, n23, n24, n25;

  BUFX10 U3 ( .A(n8), .Y(n18) );
  OAI2BB1X4TH U4 ( .A0N(n23), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI221XLTH U5 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n18), .Y(
        out[2]) );
  OAI221XLTH U6 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n18), .Y(
        out[1]) );
  INVXLTH U7 ( .A(in[4]), .Y(n22) );
  INVX2TH U8 ( .A(in[5]), .Y(n21) );
  OAI211XLTH U9 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n18), .Y(out[3]) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n23) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U13 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U15 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  XNOR2XLTH U16 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U18 ( .A(in[2]), .Y(n24) );
  INVXLTH U19 ( .A(in[6]), .Y(n20) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  OAI33X4 U21 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n21), .B2(
        n22), .Y(n8) );
endmodule


module tc_sm_120 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n19, n20, n21, n22, n23, n24, n25;

  OAI2BB1X2 U3 ( .A0N(n23), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI221XL U4 ( .A0(n20), .A1(n12), .B0(out[4]), .B1(n25), .C0(n19), .Y(out[1]) );
  BUFX8 U5 ( .A(n8), .Y(n19) );
  OAI211XL U6 ( .A0(out[4]), .A1(n23), .B0(n7), .C0(n19), .Y(out[3]) );
  BUFX2TH U7 ( .A(in[6]), .Y(out[4]) );
  CLKINVX2TH U8 ( .A(in[6]), .Y(n20) );
  OAI21XLTH U9 ( .A0(n9), .A1(n23), .B0(out[4]), .Y(n7) );
  CLKINVX1TH U10 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U12 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U14 ( .A(n24), .B(n11), .Y(n10) );
  INVXLTH U15 ( .A(in[2]), .Y(n24) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI221XLTH U17 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n19), .Y(
        out[2]) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n19), .Y(out[0]) );
  OAI33X4 U19 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n21), .B2(
        n22), .Y(n8) );
  INVXL U20 ( .A(in[5]), .Y(n21) );
  INVXL U21 ( .A(in[4]), .Y(n22) );
endmodule


module total_3_test_17 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n68, n69, w5_4_, n6, n8, n9, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_123 sm_tc_1 ( .out(a1), .in({n6, a[3:0]}) );
  sm_tc_122 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_121 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_120 sm_tc_4 ( .out(in1), .in(in) );
  add_30 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_123 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_122 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_121 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_120 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n54), .CK(clk), .RN(n8), 
        .Q(up1[3]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n59), .CK(clk), .RN(n8), 
        .Q(up3[4]) );
  SDFFRQXLTH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n50), .CK(clk), .RN(rst), 
        .Q(n69) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n55), .CK(clk), .RN(n8), .Q(
        up1[0]) );
  SDFFRQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n57), .CK(clk), .RN(n8), 
        .Q(up1[4]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n51), .CK(clk), .RN(n9), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n57), .CK(clk), .RN(n8), 
        .Q(up3[0]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n58), .CK(clk), .RN(n8), 
        .Q(up3[1]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n50), .CK(clk), .RN(n8), 
        .Q(n68) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n60), .CK(clk), .RN(n8), 
        .Q(up2[0]) );
  BUFX6 U3 ( .A(a[4]), .Y(n6) );
  BUFX3TH U4 ( .A(rst), .Y(n8) );
  CLKBUFX1TH U6 ( .A(rst), .Y(n9) );
  SDFFRX4 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n54), .CK(clk), .RN(n8), 
        .Q(up2[2]) );
  SDFFRX4 h_reg ( .D(w5_4_), .SI(test_si), .SE(n55), .CK(clk), .RN(n9), .Q(h)
         );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n51), .CK(clk), .RN(n9), 
        .Q(up1[2]) );
  SDFFRHQX8 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n60), .CK(clk), .RN(n8), 
        .Q(up1[1]) );
  SDFFRHQX8 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n58), .CK(clk), .RN(n8), 
        .Q(up3[2]) );
  SDFFRHQX8 up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n59), .CK(clk), .RN(n8), 
        .Q(up3[3]) );
  DLY1X1TH U38 ( .A(n69), .Y(up2[1]) );
  INVXLTH U39 ( .A(n53), .Y(n50) );
  INVXLTH U40 ( .A(n52), .Y(n51) );
  DLY1X1TH U41 ( .A(n56), .Y(n52) );
  DLY1X1TH U42 ( .A(n56), .Y(n53) );
  INVXLTH U43 ( .A(n53), .Y(n54) );
  INVXLTH U44 ( .A(n52), .Y(n55) );
  INVXLTH U45 ( .A(test_se), .Y(n56) );
  INVXLTH U46 ( .A(n53), .Y(n57) );
  INVXLTH U47 ( .A(n52), .Y(n58) );
  INVXLTH U48 ( .A(n53), .Y(n59) );
  INVXLTH U49 ( .A(n52), .Y(n60) );
  DLY1X1TH U50 ( .A(n68), .Y(up2[3]) );
endmodule


module sm_tc_119 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n28, n29, n30, n34, n35, n38;

  INVX4 U2 ( .A(in[4]), .Y(n35) );
  XNOR2X2 U3 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI22X1TH U4 ( .A0(in[4]), .A1(n34), .B0(n35), .B1(n5), .Y(out[2]) );
  AOI31X1 U5 ( .A0(n3), .A1(n4), .A2(n5), .B0(n35), .Y(out[4]) );
  OAI2BB2XL U6 ( .B0(n35), .B1(n4), .A0N(in[3]), .A1N(n35), .Y(out[3]) );
  CLKBUFX2TH U7 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U8 ( .A(out[4]), .Y(out[6]) );
  NAND2XLTH U9 ( .A(n8), .B(n34), .Y(n7) );
  NAND2X2TH U10 ( .A(n34), .B(n8), .Y(n29) );
  INVX2 U11 ( .A(in[2]), .Y(n34) );
  NOR2X6TH U12 ( .A(in[1]), .B(in[0]), .Y(n8) );
  NAND2X4 U13 ( .A(n29), .B(n30), .Y(n5) );
  AO21XL U14 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2X4TH U15 ( .B0(n35), .B1(n6), .A0N(in[1]), .A1N(n35), .Y(out[1]) );
  NAND2X3TH U16 ( .A(n38), .B(n28), .Y(n30) );
  INVXLTH U17 ( .A(n8), .Y(n28) );
  NOR2BXLTH U18 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKBUFX1TH U19 ( .A(out[4]), .Y(out[5]) );
  CLKINVX40 U20 ( .A(n34), .Y(n38) );
endmodule


module sm_tc_118 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n4, n5, n6, n7, n26, n29, n30, n33, n34, n35, n36, n37;

  OAI2BB2X2 U3 ( .B0(n29), .B1(n5), .A0N(in[1]), .A1N(n29), .Y(out[1]) );
  INVX2TH U6 ( .A(in[2]), .Y(n30) );
  INVX2TH U7 ( .A(in[4]), .Y(n29) );
  OAI2BB2X2TH U8 ( .B0(n29), .B1(n37), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  AO21X2TH U9 ( .A0(in[0]), .A1(in[1]), .B0(n7), .Y(n5) );
  AOI31X4TH U10 ( .A0(n6), .A1(n37), .A2(n4), .B0(n29), .Y(out[4]) );
  OAI22X2 U12 ( .A0(in[4]), .A1(n34), .B0(n29), .B1(n4), .Y(out[2]) );
  INVXLTH U13 ( .A(n26), .Y(out[6]) );
  INVXLTH U14 ( .A(out[4]), .Y(n26) );
  INVXLTH U15 ( .A(n26), .Y(out[5]) );
  NOR2BXLTH U16 ( .AN(n5), .B(in[0]), .Y(n6) );
  CLKBUFX2TH U17 ( .A(in[0]), .Y(out[0]) );
  XOR2X1 U2 ( .A(n34), .B(n35), .Y(n4) );
  CLKINVX40 U4 ( .A(n30), .Y(n33) );
  CLKINVX40 U5 ( .A(n33), .Y(n34) );
  OR2X8 U11 ( .A(in[1]), .B(in[0]), .Y(n35) );
  CLKINVX40 U18 ( .A(n35), .Y(n7) );
  XOR2X1 U19 ( .A(n36), .B(in[3]), .Y(n37) );
  CLKAND2X12 U20 ( .A(n7), .B(n34), .Y(n36) );
endmodule


module sm_tc_117 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n22, n24, n25, n27, n28;

  AO21XL U3 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  INVX4 U4 ( .A(n22), .Y(out[0]) );
  XNOR2X2 U5 ( .A(n25), .B(n8), .Y(n5) );
  AOI31X2TH U6 ( .A0(n3), .A1(n4), .A2(n5), .B0(n24), .Y(out[4]) );
  INVX2 U7 ( .A(in[4]), .Y(n24) );
  INVX2 U8 ( .A(in[2]), .Y(n25) );
  OAI2BB2X1TH U9 ( .B0(n24), .B1(n6), .A0N(in[1]), .A1N(n24), .Y(out[1]) );
  OAI22XL U10 ( .A0(in[4]), .A1(n25), .B0(n24), .B1(n5), .Y(out[2]) );
  OAI2BB2XLTH U11 ( .B0(n24), .B1(n4), .A0N(n27), .A1N(n24), .Y(out[3]) );
  NOR2X8 U13 ( .A(in[1]), .B(out[0]), .Y(n8) );
  NOR2BXLTH U14 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[6]) );
  INVX2TH U17 ( .A(in[0]), .Y(n22) );
  CLKBUFX40 U2 ( .A(in[3]), .Y(n27) );
  XOR2X1 U12 ( .A(n28), .B(n27), .Y(n4) );
  CLKAND2X12 U18 ( .A(n8), .B(n25), .Y(n28) );
endmodule


module sm_tc_116 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n18, n19, n20, n22, n25, n26;

  NOR2X4TH U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  AOI31X2TH U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n26), .Y(out[4]) );
  NAND2X1TH U4 ( .A(n8), .B(n25), .Y(n7) );
  INVXLTH U5 ( .A(n7), .Y(n17) );
  OAI2BB2X1TH U6 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  OAI2BB2X2TH U7 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n26), .Y(out[1]) );
  CLKBUFX1TH U8 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U9 ( .A(n22), .Y(out[6]) );
  OAI22X1TH U10 ( .A0(in[4]), .A1(n25), .B0(n26), .B1(n5), .Y(out[2]) );
  CLKNAND2X4 U11 ( .A(n7), .B(in[3]), .Y(n19) );
  NAND2X8 U12 ( .A(n17), .B(n18), .Y(n20) );
  NAND2X8 U13 ( .A(n19), .B(n20), .Y(n4) );
  INVXLTH U14 ( .A(in[3]), .Y(n18) );
  CLKINVX1TH U15 ( .A(in[2]), .Y(n25) );
  CLKINVX2TH U16 ( .A(in[4]), .Y(n26) );
  INVXLTH U17 ( .A(out[4]), .Y(n22) );
  NOR2BXLTH U18 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U19 ( .A(n22), .Y(out[5]) );
  XNOR2X1TH U20 ( .A(n25), .B(n8), .Y(n5) );
  AO21XLTH U21 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_29_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n4, n5, n6, n7, n8;
  wire   [6:2] carry;

  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n6), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2X1TH U1 ( .A(n4), .B(n5), .Y(SUM[0]) );
  NAND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n4) );
  NAND2XLTH U3 ( .A(n7), .B(n8), .Y(n5) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n6) );
  INVXLTH U5 ( .A(A[0]), .Y(n8) );
  INVXLTH U6 ( .A(B[0]), .Y(n7) );
endmodule


module add_29_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   carry_2_, n1;
  wire   [6:3] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry_2_), .S(SUM[1]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKAND2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_29_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_29_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_29_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_1 ( .A(B[1]), .B(n1), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X2 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_29_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_2 ( .A(carry[2]), .B(B[2]), .CI(A[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_29 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n16, n17, n18, n19, n20, n21, n22;

  add_29_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n20, n22, 
        temp1_1_, n19}), .B(in2), .SUM(out3) );
  add_29_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_29_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n20, n22, 
        temp1_1_, n19}), .B({n17, in3[5:4], n16, in3[2], n18, in3[0]}), .SUM(
        out2) );
  add_29_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n20, n22, 
        temp1_1_, n19}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_29_DW01_add_4 add_30 ( .A(in2), .B({n17, in3[5:4], n21, in3[2], n18, 
        in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_29_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX1TH U1 ( .A(n21), .Y(n16) );
  CLKBUFX1TH U2 ( .A(in3[6]), .Y(n17) );
  CLKBUFX40 U3 ( .A(in3[1]), .Y(n18) );
  CLKBUFX40 U4 ( .A(temp1_0_), .Y(n19) );
  CLKBUFX40 U5 ( .A(temp1_3_), .Y(n20) );
  CLKBUFX40 U6 ( .A(in3[3]), .Y(n21) );
  CLKBUFX40 U13 ( .A(temp1_2_), .Y(n22) );
endmodule


module tc_sm_119 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  BUFX2 U3 ( .A(in[6]), .Y(out[4]) );
  NOR3X1TH U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U5 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U6 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U7 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U8 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n28) );
  INVXLTH U12 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n29) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_118 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n16, n17, n18, n19, n20, n21;

  OAI211XL U3 ( .A0(in[6]), .A1(n19), .B0(n7), .C0(n14), .Y(out[3]) );
  BUFX10 U4 ( .A(n8), .Y(n14) );
  OAI221X1 U5 ( .A0(n16), .A1(n10), .B0(in[6]), .B1(n20), .C0(n14), .Y(out[2])
         );
  OAI33X4 U6 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n17), .B2(n18), .Y(n8) );
  OAI2BB1X4 U7 ( .A0N(n19), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI221X1TH U8 ( .A0(n16), .A1(n12), .B0(in[6]), .B1(n21), .C0(n14), .Y(
        out[1]) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n19) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U11 ( .A(n20), .B(n11), .Y(n10) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U13 ( .A(in[6]), .Y(n16) );
  OAI21XLTH U14 ( .A0(n9), .A1(n19), .B0(in[6]), .Y(n7) );
  INVX2 U15 ( .A(in[5]), .Y(n17) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U17 ( .A(in[2]), .Y(n20) );
  INVXLTH U18 ( .A(in[1]), .Y(n21) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n14), .Y(out[0]) );
  INVXL U21 ( .A(in[4]), .Y(n18) );
endmodule


module tc_sm_117 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n17, n18, n19, n20, n21, n22, n24, n25,
         n26, n27, n28;

  CLKINVX6TH U3 ( .A(n19), .Y(n8) );
  OAI221X1TH U4 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n28), .C0(n8), .Y(out[1]) );
  INVXLTH U5 ( .A(in[6]), .Y(n24) );
  AOI21BX1TH U6 ( .A0(n26), .A1(n9), .B0N(in[6]), .Y(n22) );
  NAND3XLTH U7 ( .A(n17), .B(n18), .C(n8), .Y(out[2]) );
  OR2XLTH U8 ( .A(n24), .B(n10), .Y(n17) );
  AOI33X4 U9 ( .A0(n25), .A1(n20), .A2(n21), .B0(n22), .B1(in[5]), .B2(in[4]), 
        .Y(n19) );
  OR2XLTH U10 ( .A(in[6]), .B(n27), .Y(n18) );
  INVXLTH U11 ( .A(in[6]), .Y(n20) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n26) );
  INVXLTH U14 ( .A(in[4]), .Y(n25) );
  INVXLTH U15 ( .A(in[5]), .Y(n21) );
  OAI211XLTH U16 ( .A0(in[6]), .A1(n26), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI21XLTH U17 ( .A0(n9), .A1(n26), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U18 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  XNOR2XLTH U20 ( .A(n27), .B(n11), .Y(n10) );
  NOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U22 ( .A(in[2]), .Y(n27) );
  INVXLTH U23 ( .A(in[1]), .Y(n28) );
  XNOR2XLTH U24 ( .A(in[0]), .B(in[1]), .Y(n12) );
endmodule


module tc_sm_116 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n22, n23, n24, n26, n27, n28,
         n29;

  INVXLTH U3 ( .A(in[5]), .Y(n20) );
  OAI221XL U4 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1])
         );
  OAI221XL U6 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2])
         );
  INVXLTH U7 ( .A(in[6]), .Y(n19) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n22) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U10 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U11 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI21XLTH U13 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  INVXLTH U14 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U16 ( .A(in[2]), .Y(n23) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211XLTH U18 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  AOI33X4 U5 ( .A0(n27), .A1(n28), .A2(n20), .B0(n29), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U19 ( .A(n26), .Y(n8) );
  CLKINVX40 U20 ( .A(in[4]), .Y(n27) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n28) );
  AOI21BX4 U22 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n29) );
endmodule


module total_3_test_18 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n60, n61, w5_4_, n5, n6, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_119 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_118 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_117 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_116 sm_tc_4 ( .out(in1), .in(in) );
  add_29 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_119 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_118 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_117 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_116 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(n61) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n58), .CK(clk), .RN(n6), 
        .Q(up2[4]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n53), .CK(clk), .RN(n6), .Q(
        h) );
  SDFFRQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n56), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up2[1]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n58), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  SDFFRQX2TH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n56), .CK(clk), .RN(n5), 
        .Q(up1[2]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n52), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRQXL up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n53), .CK(clk), .RN(n5), 
        .Q(up1[3]) );
  SDFFRQX1TH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n57), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRQXLTH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n55), .CK(clk), .RN(n6), .Q(
        n60) );
  SDFFRQX4 up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n52), .CK(clk), .RN(n5), 
        .Q(up3[4]) );
  SDFFRQX1TH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up3[3]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n6) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n5) );
  SDFFRX4 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up2[2]) );
  SDFFRHQX8 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n57), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  SDFFRHQX8 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n55), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  DLY1X1TH U37 ( .A(n61), .Y(up2[0]) );
  DLY1X1TH U38 ( .A(n60), .Y(up1[0]) );
  INVXLTH U39 ( .A(n50), .Y(n48) );
  INVXLTH U40 ( .A(n51), .Y(n49) );
  DLY1X1TH U41 ( .A(n54), .Y(n50) );
  DLY1X1TH U42 ( .A(n54), .Y(n51) );
  INVXLTH U43 ( .A(n51), .Y(n52) );
  INVXLTH U44 ( .A(n50), .Y(n53) );
  INVXLTH U45 ( .A(test_se), .Y(n54) );
  INVXLTH U46 ( .A(n51), .Y(n55) );
  INVXLTH U47 ( .A(n50), .Y(n56) );
  INVXLTH U48 ( .A(n51), .Y(n57) );
  INVXLTH U49 ( .A(n50), .Y(n58) );
endmodule


module sm_tc_115 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n24, n25, n28, n29, n30;

  INVX2 U2 ( .A(in[2]), .Y(n25) );
  NOR2X4 U3 ( .A(n30), .B(in[0]), .Y(n8) );
  AO21X2 U4 ( .A0(in[0]), .A1(n30), .B0(n8), .Y(n6) );
  OAI2BB2X2 U5 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  INVX3 U6 ( .A(in[4]), .Y(n24) );
  CLKBUFX1TH U7 ( .A(out[4]), .Y(out[6]) );
  AOI31X2TH U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n29), .Y(out[4]) );
  OAI2BB2X4TH U9 ( .B0(n29), .B1(n6), .A0N(n30), .A1N(n29), .Y(out[1]) );
  OAI22XL U10 ( .A0(in[4]), .A1(n25), .B0(n29), .B1(n5), .Y(out[2]) );
  XNOR2X1 U11 ( .A(n25), .B(n8), .Y(n5) );
  CLKBUFX1TH U12 ( .A(in[0]), .Y(out[0]) );
  XNOR2X2 U13 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U14 ( .A(n8), .B(n25), .Y(n7) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  CLKINVX40 U17 ( .A(n24), .Y(n28) );
  CLKINVX40 U18 ( .A(n28), .Y(n29) );
  CLKBUFX40 U19 ( .A(in[1]), .Y(n30) );
endmodule


module sm_tc_114 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n28, n29, n31;

  INVX2 U2 ( .A(in[4]), .Y(n29) );
  OAI22X1 U3 ( .A0(in[4]), .A1(n28), .B0(n29), .B1(n5), .Y(out[2]) );
  OAI2BB2X1TH U5 ( .B0(n29), .B1(n6), .A0N(in[1]), .A1N(n29), .Y(out[1]) );
  AOI31X2TH U6 ( .A0(n3), .A1(n4), .A2(n5), .B0(n29), .Y(out[6]) );
  OAI2BB2XL U7 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  NOR2BXLTH U8 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVX1TH U9 ( .A(in[2]), .Y(n28) );
  CLKBUFX1TH U10 ( .A(out[6]), .Y(out[4]) );
  XNOR2X1TH U11 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX1TH U12 ( .A(out[6]), .Y(out[5]) );
  NAND2XLTH U13 ( .A(n8), .B(n28), .Y(n7) );
  XNOR2X1TH U14 ( .A(n28), .B(n8), .Y(n5) );
  BUFX2TH U15 ( .A(in[0]), .Y(out[0]) );
  AO21XLTH U16 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OR2X8 U4 ( .A(in[1]), .B(in[0]), .Y(n31) );
  CLKINVX40 U17 ( .A(n31), .Y(n8) );
endmodule


module sm_tc_113 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n35, n3, n5, n6, n7, n8, n21, n22, n26, n27, n29, n30, n31, n32, n33;

  OAI2BB2X2 U5 ( .B0(n32), .B1(n6), .A0N(n29), .A1N(n32), .Y(out[1]) );
  INVX1TH U2 ( .A(in[2]), .Y(n27) );
  AOI31X2TH U3 ( .A0(n3), .A1(n30), .A2(n21), .B0(n32), .Y(n35) );
  BUFX6 U4 ( .A(n5), .Y(n21) );
  XNOR2XL U6 ( .A(n27), .B(n8), .Y(n5) );
  BUFX3 U7 ( .A(in[4]), .Y(n22) );
  CLKNAND2X2 U9 ( .A(n8), .B(n27), .Y(n7) );
  INVX2TH U10 ( .A(n22), .Y(n26) );
  AO21XL U11 ( .A0(in[0]), .A1(n29), .B0(n8), .Y(n6) );
  OAI22X4TH U12 ( .A0(n22), .A1(n27), .B0(n32), .B1(n21), .Y(out[2]) );
  OAI2BB2X1TH U13 ( .B0(n32), .B1(n30), .A0N(in[3]), .A1N(n32), .Y(out[3]) );
  NOR2X2 U14 ( .A(n29), .B(in[0]), .Y(n8) );
  CLKBUFX1TH U15 ( .A(out[6]), .Y(out[4]) );
  CLKBUFX1TH U16 ( .A(out[6]), .Y(out[5]) );
  BUFX2TH U17 ( .A(in[0]), .Y(out[0]) );
  NOR2BXLTH U18 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX40 U8 ( .A(in[1]), .Y(n29) );
  XNOR2X1 U19 ( .A(n7), .B(in[3]), .Y(n30) );
  CLKINVX40 U20 ( .A(n26), .Y(n31) );
  CLKINVX40 U21 ( .A(n31), .Y(n32) );
  CLKINVX40 U22 ( .A(n35), .Y(n33) );
  CLKINVX40 U23 ( .A(n33), .Y(out[6]) );
endmodule


module sm_tc_112 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  OAI2BB2X2 U2 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  XNOR2X1TH U3 ( .A(n7), .B(in[3]), .Y(n4) );
  AOI31X2TH U4 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  OAI2BB2X2TH U5 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U6 ( .A(in[0]), .Y(out[0]) );
  AO21XLTH U7 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI22X1TH U8 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  NOR2X4TH U9 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX2TH U10 ( .A(in[4]), .Y(n22) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n21) );
  INVXLTH U12 ( .A(out[4]), .Y(n18) );
  CLKINVX1TH U13 ( .A(n18), .Y(out[5]) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U15 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U16 ( .A(n21), .B(n8), .Y(n5) );
  NAND2XLTH U17 ( .A(n8), .B(n21), .Y(n7) );
endmodule


module add_28_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_28_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18;
  wire   [6:2] carry;

  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX4TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3XL U1 ( .A(A[3]), .B(carry[3]), .C(B[3]), .Y(SUM[3]) );
  NAND2X2 U2 ( .A(A[3]), .B(carry[3]), .Y(n10) );
  NAND2XL U3 ( .A(A[3]), .B(B[3]), .Y(n11) );
  NAND2X2 U4 ( .A(carry[3]), .B(B[3]), .Y(n12) );
  NAND3X2 U5 ( .A(n10), .B(n11), .C(n12), .Y(carry[4]) );
  NAND2XLTH U7 ( .A(A[1]), .B(n1), .Y(n7) );
  INVXLTH U8 ( .A(n6), .Y(n15) );
  CLKNAND2X2TH U9 ( .A(n15), .B(A[1]), .Y(n5) );
  NAND2XLTH U10 ( .A(n6), .B(n14), .Y(n4) );
  NAND3X2TH U11 ( .A(n7), .B(n8), .C(n9), .Y(carry[2]) );
  NAND2XLTH U12 ( .A(n1), .B(B[1]), .Y(n9) );
  CLKXOR2X1TH U13 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X1TH U14 ( .A(B[0]), .B(A[0]), .Y(n1) );
  NAND2XLTH U15 ( .A(A[1]), .B(B[1]), .Y(n8) );
  INVXLTH U16 ( .A(A[1]), .Y(n14) );
  CLKXOR2X4 U17 ( .A(B[6]), .B(A[6]), .Y(n13) );
  CLKXOR2X12 U18 ( .A(n13), .B(carry[6]), .Y(SUM[6]) );
  AND2X8 U6 ( .A(n4), .B(n5), .Y(n16) );
  CLKINVX40 U19 ( .A(n16), .Y(SUM[1]) );
  DLY1X1TH U20 ( .A(n18), .Y(n17) );
  XNOR2X1 U21 ( .A(B[1]), .B(n1), .Y(n18) );
  CLKINVX40 U22 ( .A(n17), .Y(n6) );
endmodule


module add_28_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_28_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(n2), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKINVX40 U4 ( .A(A[6]), .Y(n2) );
endmodule


module add_28_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  CLKXOR2X2TH U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFHXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(carry[3]), .CI(B[3]), .CO(carry[4]), .S(SUM[3])
         );
  CLKXOR2X2TH U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XLTH U4 ( .A(B[6]), .B(A[6]), .Y(n2) );
endmodule


module add_28_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX2 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR2X3TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_28 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n18, n19, n20, n21, n22;

  add_28_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, n21, temp1_3_, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in2[6:3], n19, n18, in2[0]}), .SUM(out3) );
  add_28_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_28_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, n20, temp1_3_, temp1_2_, 
        temp1_1_, temp1_0_}), .B(in3), .SUM(out2) );
  add_28_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, n22, temp1_3_, temp1_2_, 
        temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_28_DW01_add_4 add_30 ( .A({in2[6:3], n19, n18, in2[0]}), .B(in3), .SUM({
        temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_})
         );
  add_28_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX2TH U1 ( .A(in2[2]), .Y(n19) );
  BUFX2TH U2 ( .A(in2[1]), .Y(n18) );
  CLKBUFX1TH U3 ( .A(n21), .Y(n20) );
  CLKBUFX40 U4 ( .A(temp1_4_), .Y(n21) );
  CLKBUFX1TH U5 ( .A(n21), .Y(n22) );
endmodule


module tc_sm_115 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n23, n25, n26, n27, n28, n29, n30;

  CLKBUFX2TH U3 ( .A(in[6]), .Y(n23) );
  NOR3X1TH U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U5 ( .A(in[1]), .Y(n30) );
  XNOR2XLTH U6 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U7 ( .A(in[2]), .Y(n29) );
  XNOR2XLTH U8 ( .A(n29), .B(n11), .Y(n10) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(n23), .A2(in[5]), .B0(n13), .B1(n26), .B2(
        n27), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n27) );
  INVXLTH U12 ( .A(in[5]), .Y(n26) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n28) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U15 ( .A(n23), .Y(n25) );
  OAI221XLTH U16 ( .A0(n25), .A1(n12), .B0(n23), .B1(n30), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U17 ( .A0(n25), .A1(n10), .B0(n23), .B1(n29), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U18 ( .A0(n9), .A1(n28), .B0(n23), .Y(n7) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211XLTH U20 ( .A0(n23), .A1(n28), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U21 ( .A0N(n28), .A1N(n9), .B0(n23), .Y(n13) );
endmodule


module tc_sm_114 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n20, n22, n23, n24, n25, n26, n27;

  BUFX10 U3 ( .A(n8), .Y(n20) );
  OAI221X2 U4 ( .A0(n22), .A1(n10), .B0(in[6]), .B1(n26), .C0(n20), .Y(out[2])
         );
  OAI2BB1X4 U5 ( .A0N(n25), .A1N(n9), .B0(in[6]), .Y(n13) );
  NAND2BX1TH U6 ( .AN(in[0]), .B(n20), .Y(out[0]) );
  OAI221X2 U7 ( .A0(n22), .A1(n12), .B0(in[6]), .B1(n27), .C0(n20), .Y(out[1])
         );
  OAI211X2 U8 ( .A0(in[6]), .A1(n25), .B0(n7), .C0(n20), .Y(out[3]) );
  INVXLTH U9 ( .A(in[6]), .Y(n22) );
  INVX2TH U10 ( .A(in[4]), .Y(n24) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n25) );
  INVXLTH U12 ( .A(in[1]), .Y(n27) );
  XNOR2XLTH U13 ( .A(n26), .B(n11), .Y(n10) );
  INVXLTH U14 ( .A(in[2]), .Y(n26) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U16 ( .A0(n9), .A1(n25), .B0(in[6]), .Y(n7) );
  INVX2 U17 ( .A(in[5]), .Y(n23) );
  XNOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n11) );
  NOR3X1TH U20 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  OAI33X4 U21 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n23), .B2(
        n24), .Y(n8) );
endmodule


module tc_sm_113 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n20, n21, n22, n23, n24, n25,
         n27;

  BUFX5 U3 ( .A(n8), .Y(n18) );
  OAI2BB1X2TH U4 ( .A0N(n23), .A1N(n9), .B0(n27), .Y(n13) );
  INVXLTH U5 ( .A(n27), .Y(n20) );
  CLKINVX1TH U6 ( .A(in[3]), .Y(n23) );
  OAI221XLTH U7 ( .A0(n20), .A1(n10), .B0(n27), .B1(n24), .C0(n18), .Y(out[2])
         );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U9 ( .A(n27), .Y(out[4]) );
  XNOR2XLTH U10 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U12 ( .A(in[2]), .Y(n24) );
  OAI21XLTH U13 ( .A0(n9), .A1(n23), .B0(n27), .Y(n7) );
  INVXLTH U14 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI221XLTH U16 ( .A0(n20), .A1(n12), .B0(n27), .B1(n25), .C0(n18), .Y(out[1]) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  OAI211XLTH U18 ( .A0(n27), .A1(n23), .B0(n7), .C0(n18), .Y(out[3]) );
  OAI33X4 U19 ( .A0(in[4]), .A1(n27), .A2(in[5]), .B0(n13), .B1(n21), .B2(n22), 
        .Y(n8) );
  INVXL U20 ( .A(in[5]), .Y(n21) );
  INVXL U21 ( .A(in[4]), .Y(n22) );
  CLKBUFX40 U22 ( .A(in[6]), .Y(n27) );
endmodule


module tc_sm_112 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n20, n21, n22, n23, n24, n25;

  OAI211X1 U3 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n18), .Y(out[3]) );
  BUFX10 U4 ( .A(n8), .Y(n18) );
  OAI221XL U5 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n18), .Y(out[1])
         );
  OAI2BB1X4 U6 ( .A0N(n23), .A1N(n9), .B0(in[6]), .Y(n13) );
  INVXLTH U7 ( .A(in[5]), .Y(n21) );
  OAI221X1TH U8 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n18), .Y(
        out[2]) );
  INVXLTH U9 ( .A(in[6]), .Y(n20) );
  CLKINVX1TH U10 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U12 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI21XLTH U14 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  INVXLTH U15 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U18 ( .A(in[2]), .Y(n24) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  OAI33X4 U20 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n21), .B2(
        n22), .Y(n8) );
  INVXL U21 ( .A(in[4]), .Y(n22) );
endmodule


module total_3_test_19 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n61, w5_4_, n6, n7, n8, n9, n44, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_115 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_114 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_113 sm_tc_3 ( .out(c1), .in({c[4:1], n7}) );
  sm_tc_112 sm_tc_4 ( .out(in1), .in(in) );
  add_28 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3({c1[6:2], n44, c1[0]}), .in(in1) );
  tc_sm_115 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_114 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_113 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_112 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n46), .CK(clk), .RN(n9), 
        .Q(up3[3]) );
  SDFFRQXLTH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n56), .CK(clk), .RN(n9), 
        .Q(up1[4]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n47), .CK(clk), .RN(n8), 
        .Q(up3[2]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n50), .CK(clk), .RN(n9), .Q(
        h) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n51), .CK(clk), .RN(n8), 
        .Q(up1[3]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n56), .CK(clk), .RN(n8), 
        .Q(n61) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n54), .CK(clk), .RN(n8), 
        .Q(up3[4]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n53), .CK(clk), .RN(n8), 
        .Q(up3[0]) );
  SDFFRQXLTH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n47), .CK(clk), .RN(n8), 
        .Q(up1[1]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n54), .CK(clk), .RN(n8), 
        .Q(up2[0]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n55), .CK(clk), .RN(n8), 
        .Q(up3[1]) );
  SDFFRQX2 up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n53), .CK(clk), .RN(n8), 
        .Q(up2[4]) );
  SDFFRQX1 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n46), .CK(clk), .RN(n8), 
        .Q(up2[1]) );
  SDFFRQX4 up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n51), .CK(clk), .RN(n8), .Q(
        up1[0]) );
  INVX2TH U3 ( .A(c[0]), .Y(n6) );
  INVX1TH U4 ( .A(n6), .Y(n7) );
  CLKBUFX1TH U5 ( .A(rst), .Y(n9) );
  CLKBUFX4TH U6 ( .A(rst), .Y(n8) );
  SDFFRX4 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n50), .CK(clk), .RN(n8), 
        .Q(up2[2]) );
  SDFFRX4 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n55), .CK(clk), .RN(n8), 
        .Q(up2[3]) );
  CLKBUFX40 U39 ( .A(c1[1]), .Y(n44) );
  DLY1X1TH U40 ( .A(n61), .Y(up1[2]) );
  INVXLTH U41 ( .A(n49), .Y(n46) );
  INVXLTH U42 ( .A(n48), .Y(n47) );
  DLY1X1TH U43 ( .A(n52), .Y(n48) );
  DLY1X1TH U44 ( .A(n52), .Y(n49) );
  INVXLTH U45 ( .A(n49), .Y(n50) );
  INVXLTH U46 ( .A(n48), .Y(n51) );
  INVXLTH U47 ( .A(test_se), .Y(n52) );
  INVXLTH U48 ( .A(n49), .Y(n53) );
  INVXLTH U49 ( .A(n48), .Y(n54) );
  INVXLTH U50 ( .A(n49), .Y(n55) );
  INVXLTH U51 ( .A(n48), .Y(n56) );
endmodule


module sm_tc_111 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n19, n20, n21, n25, n26, n28, n29;

  OAI22X1 U2 ( .A0(in[4]), .A1(n26), .B0(n25), .B1(n5), .Y(out[2]) );
  NOR2X6 U3 ( .A(n29), .B(in[0]), .Y(n8) );
  CLKBUFX1TH U4 ( .A(out[6]), .Y(out[5]) );
  AOI31X2 U5 ( .A0(n3), .A1(n4), .A2(n5), .B0(n25), .Y(out[6]) );
  CLKNAND2X12 U6 ( .A(n26), .B(n8), .Y(n20) );
  AO21X2 U7 ( .A0(in[0]), .A1(n29), .B0(n8), .Y(n6) );
  NAND2XLTH U8 ( .A(n8), .B(n26), .Y(n7) );
  CLKNAND2X2 U9 ( .A(n20), .B(n21), .Y(n5) );
  INVX2 U10 ( .A(in[2]), .Y(n26) );
  INVX4TH U11 ( .A(in[4]), .Y(n25) );
  CLKINVX4 U12 ( .A(n8), .Y(n19) );
  BUFX2TH U13 ( .A(in[0]), .Y(out[0]) );
  NAND2X2 U14 ( .A(n28), .B(n19), .Y(n21) );
  OAI2BB2X4TH U15 ( .B0(n25), .B1(n6), .A0N(n29), .A1N(n25), .Y(out[1]) );
  XNOR2X4 U16 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX1TH U17 ( .A(out[6]), .Y(out[4]) );
  OAI2BB2XLTH U18 ( .B0(n25), .B1(n4), .A0N(in[3]), .A1N(n25), .Y(out[3]) );
  NOR2BXLTH U19 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX40 U20 ( .A(n26), .Y(n28) );
  CLKBUFX40 U21 ( .A(in[1]), .Y(n29) );
endmodule


module sm_tc_110 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n26, n27, n30, n31, n32;

  OAI22X2 U2 ( .A0(in[4]), .A1(n30), .B0(n26), .B1(n5), .Y(out[2]) );
  OAI2BB2X2 U4 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  CLKBUFX1TH U5 ( .A(out[4]), .Y(out[6]) );
  NAND2XLTH U6 ( .A(n8), .B(n30), .Y(n7) );
  INVX1TH U7 ( .A(in[2]), .Y(n27) );
  INVX2TH U8 ( .A(in[4]), .Y(n26) );
  XNOR2X2 U9 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X2 U10 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n26), .Y(out[1]) );
  AO21XLTH U11 ( .A0(n32), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKBUFX1TH U12 ( .A(n32), .Y(out[0]) );
  AOI31X2TH U13 ( .A0(n3), .A1(n4), .A2(n5), .B0(n26), .Y(out[4]) );
  NOR2BXLTH U14 ( .AN(n6), .B(n32), .Y(n3) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  XNOR2X1TH U16 ( .A(n30), .B(n8), .Y(n5) );
  CLKBUFX40 U3 ( .A(n27), .Y(n30) );
  OR2X8 U17 ( .A(in[1]), .B(n32), .Y(n31) );
  CLKINVX40 U18 ( .A(n31), .Y(n8) );
  CLKBUFX40 U19 ( .A(in[0]), .Y(n32) );
endmodule


module sm_tc_109 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n30, n31, n34, n35, n36;

  XNOR2X1 U3 ( .A(n7), .B(in[3]), .Y(n4) );
  BUFX5TH U4 ( .A(in[0]), .Y(out[0]) );
  INVX2 U6 ( .A(in[4]), .Y(n31) );
  AOI31X2 U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n35), .Y(out[4]) );
  OAI2BB2XL U8 ( .B0(n35), .B1(n4), .A0N(in[3]), .A1N(n35), .Y(out[3]) );
  CLKINVX1TH U9 ( .A(in[2]), .Y(n30) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[5]) );
  OAI22X2 U12 ( .A0(in[4]), .A1(n30), .B0(n35), .B1(n5), .Y(out[2]) );
  NOR2BXLTH U13 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[6]) );
  NAND2XLTH U15 ( .A(n8), .B(n30), .Y(n7) );
  AO21XLTH U16 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKINVX40 U2 ( .A(n31), .Y(n34) );
  CLKINVX40 U5 ( .A(n34), .Y(n35) );
  XOR2X1 U10 ( .A(n30), .B(n36), .Y(n5) );
  AO2B2X4 U17 ( .B0(in[1]), .B1(n35), .A0(in[4]), .A1N(n6), .Y(out[1]) );
  OR2X8 U18 ( .A(in[1]), .B(out[0]), .Y(n36) );
  CLKINVX40 U19 ( .A(n36), .Y(n8) );
endmodule


module sm_tc_108 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n24, n28, n29, n31;

  NOR2X2 U2 ( .A(n24), .B(n29), .Y(out[6]) );
  NAND2X2 U3 ( .A(n8), .B(n28), .Y(n7) );
  CLKBUFX2TH U4 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1TH U5 ( .A(n7), .B(in[3]), .Y(n4) );
  NOR2X3TH U6 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKBUFX1TH U7 ( .A(n31), .Y(out[4]) );
  AND3XLTH U8 ( .A(n3), .B(n4), .C(n5), .Y(n24) );
  OAI2BB2X1TH U9 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  OAI2BB2X2TH U10 ( .B0(n29), .B1(n6), .A0N(in[1]), .A1N(n29), .Y(out[1]) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n28) );
  XNOR2X1TH U12 ( .A(n28), .B(n8), .Y(n5) );
  CLKINVX2TH U13 ( .A(in[4]), .Y(n29) );
  CLKBUFX1TH U14 ( .A(n31), .Y(out[5]) );
  OAI22X4TH U15 ( .A0(in[4]), .A1(n28), .B0(n29), .B1(n5), .Y(out[2]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X2 U18 ( .A(n24), .B(n29), .Y(n31) );
endmodule


module add_27_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_27_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7;
  wire   [6:2] carry;

  ADDFHX4TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n5), .CO(carry[2]), .S(SUM[1]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  NAND2XLTH U1 ( .A(carry[2]), .B(B[2]), .Y(n4) );
  NAND3X2TH U2 ( .A(n2), .B(n3), .C(n4), .Y(carry[3]) );
  NAND2XLTH U3 ( .A(A[2]), .B(carry[2]), .Y(n2) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n5) );
  CLKXOR2X1TH U5 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  CLKXOR2X1TH U6 ( .A(n1), .B(A[2]), .Y(SUM[2]) );
  XOR2XLTH U7 ( .A(B[2]), .B(carry[2]), .Y(n1) );
  NAND2XLTH U8 ( .A(A[2]), .B(B[2]), .Y(n3) );
  XOR3X2 U9 ( .A(A[6]), .B(n6), .C(carry[6]), .Y(n7) );
  CLKINVX40 U10 ( .A(B[6]), .Y(n6) );
  CLKINVX40 U11 ( .A(n7), .Y(SUM[6]) );
endmodule


module add_27_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3;
  wire   [6:2] carry;

  ADDFHXLTH U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X2 U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U4 ( .A(A[0]), .B(B[0]), .Y(n1) );
  XNOR2X1 U3 ( .A(n3), .B(A[6]), .Y(n2) );
  CLKINVX40 U5 ( .A(B[6]), .Y(n3) );
endmodule


module add_27_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_27_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_1 ( .A(B[1]), .B(A[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_27_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n7, n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2TH U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(n7) );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  NAND2X4TH U1 ( .A(n4), .B(n5), .Y(SUM[0]) );
  NAND2XL U2 ( .A(B[0]), .B(n3), .Y(n4) );
  CLKNAND2X4 U3 ( .A(n2), .B(A[0]), .Y(n5) );
  INVX4 U4 ( .A(B[0]), .Y(n2) );
  INVXLTH U5 ( .A(A[0]), .Y(n3) );
  AND2XLTH U6 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKBUFX40 U7 ( .A(n7), .Y(SUM[3]) );
endmodule


module add_27 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n22, n23, n24, n25, n27, n28, n29, n30, n31, n32, n33;

  add_27_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in2[6:4], n27, in2[2], n29, n33}), 
        .SUM(out3) );
  add_27_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, n32, temp2_2_, 
        temp2_1_, temp2_0_}), .B({in[6:5], n30, in[3:0]}), .SUM(out1) );
  add_27_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({n31, in3[5:4], n22, in3[2:0]}), 
        .SUM(out2) );
  add_27_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, n24, temp1_3_, temp1_2_, 
        temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, n32, temp2_2_, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_27_DW01_add_4 add_30 ( .A({in2[6:2], n29, n33}), .B({n28, in3[5:4], n22, 
        in3[2:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_27_DW01_add_5 add_29 ( .A({in[6:5], n30, in[3:0]}), .B(in1), .SUM({
        temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_})
         );
  BUFX2 U1 ( .A(in3[3]), .Y(n22) );
  INVXLTH U2 ( .A(in2[3]), .Y(n25) );
  INVXLTH U3 ( .A(temp1_4_), .Y(n23) );
  INVXLTH U4 ( .A(n23), .Y(n24) );
  INVXLTH U6 ( .A(n25), .Y(n27) );
  CLKBUFX1TH U13 ( .A(in3[6]), .Y(n28) );
  CLKBUFX40 U5 ( .A(in2[1]), .Y(n29) );
  DLY1X1TH U14 ( .A(in[4]), .Y(n30) );
  CLKBUFX1TH U15 ( .A(in3[6]), .Y(n31) );
  CLKBUFX40 U16 ( .A(temp2_3_), .Y(n32) );
  CLKBUFX40 U17 ( .A(in2[0]), .Y(n33) );
endmodule


module tc_sm_111 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31, n33;

  CLKBUFX2TH U3 ( .A(n33), .Y(out[4]) );
  NOR3X1TH U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U5 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U6 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U7 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U8 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(n33), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n28) );
  INVXLTH U12 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n29) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(n33), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(n33), .B1(n31), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(n33), .B1(n30), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(n33), .Y(n7) );
  OAI2BB1XLTH U19 ( .A0N(n29), .A1N(n9), .B0(n33), .Y(n13) );
  OAI211XLTH U20 ( .A0(n33), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  CLKBUFX40 U21 ( .A(in[6]), .Y(n33) );
endmodule


module tc_sm_110 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n29, n30, n31, n32, n34, n35;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[5]), .C0(in[4]), .Y(n11) );
  OAI211XL U3 ( .A0(in[6]), .A1(n30), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI221XL U4 ( .A0(n29), .A1(n8), .B0(in[6]), .B1(n31), .C0(n6), .Y(out[2])
         );
  CLKINVX1 U5 ( .A(in[6]), .Y(n29) );
  OAI21X1 U6 ( .A0(n7), .A1(n30), .B0(in[6]), .Y(n5) );
  AOI21X8 U9 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n6) );
  AOI2BB1X4 U10 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  XOR2XLTH U13 ( .A(in[0]), .B(n32), .Y(n10) );
  INVXLTH U14 ( .A(in[1]), .Y(n32) );
  INVXLTH U15 ( .A(in[2]), .Y(n31) );
  XOR2XLTH U16 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n9) );
  INVXLTH U18 ( .A(in[3]), .Y(n30) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  OR2X8 U8 ( .A(n29), .B(n10), .Y(n34) );
  OR2X8 U20 ( .A(in[6]), .B(n32), .Y(n35) );
  NAND3X8 U21 ( .A(n34), .B(n35), .C(n6), .Y(out[1]) );
endmodule


module tc_sm_109 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n31, n32, n34, n35, n36, n37, n38,
         n39, n41;

  BUFX8 U3 ( .A(n8), .Y(n31) );
  CLKBUFX1TH U4 ( .A(in[6]), .Y(n32) );
  BUFX2 U6 ( .A(in[6]), .Y(out[4]) );
  OAI221X2TH U7 ( .A0(n34), .A1(n10), .B0(out[4]), .B1(n38), .C0(n31), .Y(
        out[2]) );
  OAI2BB1X4TH U8 ( .A0N(n37), .A1N(n9), .B0(n32), .Y(n13) );
  OAI221X2TH U9 ( .A0(n34), .A1(n12), .B0(out[4]), .B1(n39), .C0(n31), .Y(
        out[1]) );
  INVX2TH U10 ( .A(in[5]), .Y(n35) );
  OAI33X4 U11 ( .A0(in[4]), .A1(out[4]), .A2(in[5]), .B0(n13), .B1(n36), .B2(
        n35), .Y(n8) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n37) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U14 ( .A(in[4]), .Y(n36) );
  INVXLTH U15 ( .A(in[1]), .Y(n39) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U17 ( .A(n38), .B(n11), .Y(n10) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U19 ( .A(in[2]), .Y(n38) );
  OAI21XLTH U20 ( .A0(n9), .A1(n37), .B0(out[4]), .Y(n7) );
  NAND2BXLTH U21 ( .AN(in[0]), .B(n31), .Y(out[0]) );
  INVXLTH U22 ( .A(out[4]), .Y(n34) );
  OA21X4 U5 ( .A0(out[4]), .A1(n37), .B0(n7), .Y(n41) );
  NAND2X8 U23 ( .A(n41), .B(n31), .Y(out[3]) );
endmodule


module tc_sm_108 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n23, n24, n25, n26, n27, n28,
         n30, n31, n32;

  OAI221XL U3 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n27), .C0(n8), .Y(out[2])
         );
  OR2X2 U4 ( .A(n23), .B(n12), .Y(n20) );
  OR2XLTH U5 ( .A(in[6]), .B(n28), .Y(n21) );
  NAND3XLTH U6 ( .A(n20), .B(n21), .C(n8), .Y(out[1]) );
  OAI211XLTH U7 ( .A0(in[6]), .A1(n26), .B0(n7), .C0(n8), .Y(out[3]) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n26) );
  INVXLTH U10 ( .A(in[6]), .Y(n23) );
  INVXLTH U12 ( .A(in[1]), .Y(n28) );
  XNOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U14 ( .A(n27), .B(n11), .Y(n10) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[2]), .Y(n27) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n26), .B0(in[6]), .Y(n7) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXL U21 ( .A(in[5]), .Y(n24) );
  INVXL U22 ( .A(in[4]), .Y(n25) );
  AOI33X4 U11 ( .A0(n25), .A1(n31), .A2(n24), .B0(n32), .B1(in[5]), .B2(in[4]), 
        .Y(n30) );
  CLKINVX40 U20 ( .A(n30), .Y(n8) );
  CLKINVX40 U23 ( .A(in[6]), .Y(n31) );
  AOI21BX4 U24 ( .A0(n26), .A1(n9), .B0N(in[6]), .Y(n32) );
endmodule


module total_3_test_20 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n63, w5_4_, n7, n8, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_111 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_110 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_109 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_108 sm_tc_4 ( .out(in1), .in(in) );
  add_27 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in({in1[6:5], in1[6], in1[3:0]}) );
  tc_sm_111 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_110 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_109 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_108 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n59), .CK(clk), .RN(n7), 
        .Q(n63) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n49), .CK(clk), .RN(n7), 
        .Q(up3[0]) );
  SDFFRQX1TH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n59), .CK(clk), .RN(n7), 
        .Q(up3[2]) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n50), .CK(clk), .RN(n7), 
        .Q(up2[1]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n53), .CK(clk), .RN(n7), 
        .Q(up2[0]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n58), .CK(clk), .RN(n7), .Q(
        up1[0]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n57), .CK(clk), .RN(n7), 
        .Q(up2[3]) );
  SDFFRQX2 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n58), .CK(clk), .RN(n7), 
        .Q(up3[1]) );
  SDFFRQX2 up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n57), .CK(clk), .RN(n8), 
        .Q(up3[4]) );
  SDFFRQX1 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n54), .CK(clk), .RN(n7), 
        .Q(up1[1]) );
  SDFFRQX4TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n49), .CK(clk), .RN(n7), 
        .Q(up1[4]) );
  SDFFRQX2 up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n56), .CK(clk), .RN(n8), 
        .Q(up2[4]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n8) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n7) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n53), .CK(clk), .RN(n7), 
        .Q(up1[2]) );
  SDFFRX4 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n54), .CK(clk), .RN(n7), 
        .Q(up2[2]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n50), .CK(clk), .RN(n7), 
        .Q(up1[3]) );
  SDFFRX4 h_reg ( .D(w5_4_), .SI(test_si), .SE(n56), .CK(clk), .RN(n8), .Q(h)
         );
  INVXLTH U37 ( .A(n52), .Y(n49) );
  INVXLTH U38 ( .A(n51), .Y(n50) );
  DLY1X1TH U39 ( .A(n55), .Y(n51) );
  DLY1X1TH U40 ( .A(n55), .Y(n52) );
  INVXLTH U41 ( .A(n52), .Y(n53) );
  INVXLTH U42 ( .A(n51), .Y(n54) );
  INVXLTH U43 ( .A(test_se), .Y(n55) );
  INVXLTH U44 ( .A(n52), .Y(n56) );
  INVXLTH U45 ( .A(n51), .Y(n57) );
  INVXLTH U46 ( .A(n52), .Y(n58) );
  INVXLTH U47 ( .A(n51), .Y(n59) );
  DLY1X1TH U48 ( .A(n63), .Y(up3[3]) );
endmodule


module sm_tc_107 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n22, n23, n26;

  OAI2BB2X2 U5 ( .B0(n22), .B1(n6), .A0N(n26), .A1N(n22), .Y(out[1]) );
  NOR2X4TH U2 ( .A(n26), .B(in[0]), .Y(n8) );
  INVX2TH U3 ( .A(in[2]), .Y(n23) );
  XNOR2X1 U4 ( .A(n7), .B(in[3]), .Y(n4) );
  AO21X2TH U6 ( .A0(in[0]), .A1(n26), .B0(n8), .Y(n6) );
  AOI31X2TH U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  OAI22X2TH U8 ( .A0(n18), .A1(n23), .B0(n22), .B1(n5), .Y(out[2]) );
  NAND2XLTH U9 ( .A(n8), .B(n23), .Y(n7) );
  INVX4TH U10 ( .A(in[4]), .Y(n22) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  INVXLTH U12 ( .A(n22), .Y(n18) );
  XNOR2X1TH U13 ( .A(n23), .B(n8), .Y(n5) );
  CLKBUFX1TH U14 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2XLTH U16 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX40 U18 ( .A(in[1]), .Y(n26) );
endmodule


module sm_tc_106 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n24, n25, n29, n30, n33, n34, n35, n36, n37,
         n38;

  XNOR2X1 U2 ( .A(n34), .B(n8), .Y(n5) );
  NOR2X2 U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX2TH U4 ( .A(in[4]), .Y(n29) );
  OAI2BB2X2TH U5 ( .B0(n38), .B1(n6), .A0N(in[1]), .A1N(n38), .Y(out[1]) );
  NAND2X2TH U6 ( .A(n24), .B(n25), .Y(out[2]) );
  CLKBUFX2TH U7 ( .A(in[0]), .Y(out[0]) );
  OR2X1 U8 ( .A(n38), .B(n5), .Y(n25) );
  AOI31X4 U9 ( .A0(n3), .A1(n4), .A2(n5), .B0(n38), .Y(out[4]) );
  AO21XLTH U11 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKINVX1TH U12 ( .A(in[2]), .Y(n30) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U15 ( .A(out[5]), .Y(out[6]) );
  OR2XLTH U16 ( .A(in[4]), .B(n34), .Y(n24) );
  NAND2XLTH U17 ( .A(n8), .B(n34), .Y(n7) );
  NOR2BXLTH U18 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2B2X2 U10 ( .A1N(in[3]), .A0(n37), .B0(n38), .B1(n4), .Y(out[3]) );
  CLKBUFX40 U13 ( .A(n35), .Y(n33) );
  CLKBUFX40 U19 ( .A(n30), .Y(n34) );
  DLY1X1TH U20 ( .A(n36), .Y(n35) );
  XOR2X1 U21 ( .A(n7), .B(in[3]), .Y(n36) );
  CLKINVX40 U22 ( .A(n33), .Y(n4) );
  CLKINVX40 U23 ( .A(n29), .Y(n37) );
  CLKINVX40 U24 ( .A(n37), .Y(n38) );
endmodule


module sm_tc_105 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n23, n24, n27;

  NOR2X4 U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  AOI31X2TH U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n24), .Y(out[4]) );
  BUFX2 U4 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X2 U5 ( .B0(n24), .B1(n6), .A0N(in[1]), .A1N(n24), .Y(out[1]) );
  NAND2XL U6 ( .A(n8), .B(n23), .Y(n7) );
  INVX4TH U8 ( .A(n22), .Y(n24) );
  OAI22X4TH U9 ( .A0(n22), .A1(n23), .B0(n24), .B1(n5), .Y(out[2]) );
  XNOR2X1TH U10 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX2TH U11 ( .A(in[4]), .Y(n22) );
  INVX1TH U12 ( .A(in[2]), .Y(n23) );
  OAI2BB2X1TH U13 ( .B0(n24), .B1(n4), .A0N(in[3]), .A1N(n24), .Y(out[3]) );
  AO21XLTH U14 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[6]) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  XOR2X1 U7 ( .A(n23), .B(n27), .Y(n5) );
  CLKINVX40 U18 ( .A(n8), .Y(n27) );
endmodule


module sm_tc_104 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  CLKBUFX1TH U2 ( .A(in[0]), .Y(out[0]) );
  AOI31X4TH U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  OAI2BB2X1TH U4 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  XNOR2X2TH U5 ( .A(n7), .B(in[3]), .Y(n4) );
  NOR2X1TH U6 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U7 ( .A(in[2]), .Y(n21) );
  INVXLTH U8 ( .A(out[4]), .Y(n18) );
  XNOR2X1TH U9 ( .A(n21), .B(n8), .Y(n5) );
  CLKINVX2TH U10 ( .A(in[4]), .Y(n22) );
  CLKINVX1TH U11 ( .A(n18), .Y(out[5]) );
  OAI2BB2X2TH U12 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  OAI22X4TH U13 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  INVXLTH U14 ( .A(n18), .Y(out[6]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  NAND2XLTH U16 ( .A(n8), .B(n21), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_26_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(B[1]), .B(A[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3X4TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_26_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [6:2] carry;

  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  NAND3X4 U1 ( .A(n2), .B(n3), .C(n4), .Y(carry[2]) );
  NAND2XL U2 ( .A(A[1]), .B(B[1]), .Y(n3) );
  NAND2X2 U3 ( .A(carry[2]), .B(B[2]), .Y(n8) );
  NAND3X2 U4 ( .A(n10), .B(n11), .C(n12), .Y(carry[5]) );
  NAND2X2 U5 ( .A(A[4]), .B(carry[4]), .Y(n10) );
  NAND2XLTH U6 ( .A(A[1]), .B(n9), .Y(n2) );
  NAND3X4 U7 ( .A(n6), .B(n7), .C(n8), .Y(carry[3]) );
  NAND2XL U8 ( .A(carry[4]), .B(B[4]), .Y(n12) );
  CLKXOR2X1TH U9 ( .A(n1), .B(A[1]), .Y(SUM[1]) );
  AND2X1TH U10 ( .A(B[0]), .B(A[0]), .Y(n9) );
  XOR2XLTH U11 ( .A(B[1]), .B(n9), .Y(n1) );
  CLKXOR2X2TH U12 ( .A(n5), .B(A[2]), .Y(SUM[2]) );
  CLKNAND2X2TH U13 ( .A(A[2]), .B(B[2]), .Y(n7) );
  CLKXOR2X1TH U14 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2XLTH U15 ( .A(n9), .B(B[1]), .Y(n4) );
  CLKNAND2X2 U16 ( .A(A[2]), .B(carry[2]), .Y(n6) );
  NAND2XLTH U17 ( .A(A[4]), .B(B[4]), .Y(n11) );
  XOR2XLTH U18 ( .A(B[2]), .B(carry[2]), .Y(n5) );
  XOR3XL U19 ( .A(A[4]), .B(carry[4]), .C(B[4]), .Y(SUM[4]) );
endmodule


module add_26_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_26_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR2XL U1 ( .A(A[6]), .B(B[6]), .Y(n2) );
  CLKXOR2X4 U2 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  AND2XLTH U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_26_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n9, n1, n3, n4, n5, n6, n7;
  wire   [6:2] carry;

  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHX4 U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3XL U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX4TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XNOR2X4TH U1 ( .A(n6), .B(A[2]), .Y(n9) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR2X2TH U3 ( .A(carry[2]), .B(B[2]), .Y(n6) );
  CLKXOR2X1TH U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND3X2TH U5 ( .A(n3), .B(n4), .C(n5), .Y(carry[3]) );
  NAND2XLTH U6 ( .A(B[2]), .B(carry[2]), .Y(n5) );
  NAND2XLTH U7 ( .A(A[2]), .B(carry[2]), .Y(n4) );
  NAND2XLTH U8 ( .A(A[2]), .B(B[2]), .Y(n3) );
  CLKINVX40 U9 ( .A(n9), .Y(n7) );
  CLKINVX40 U10 ( .A(n7), .Y(SUM[2]) );
endmodule


module add_26_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n6, n7, n8, n9, n1;
  wire   [6:2] carry;

  ADDFX1TH U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(n8) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(n6) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(n9) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(n7) );
  ADDFX2TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKBUFX40 U3 ( .A(n7), .Y(SUM[4]) );
  CLKBUFX40 U4 ( .A(n9), .Y(SUM[1]) );
  CLKBUFX40 U5 ( .A(n6), .Y(SUM[5]) );
  CLKBUFX40 U6 ( .A(n8), .Y(SUM[3]) );
endmodule


module add_26 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   n27, temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_,
         temp2_0_, temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_,
         temp1_0_, n19, n21, n22, n23, n24, n25;

  add_26_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in2[6:5], n21, n24, n25, in2[1:0]}), .SUM({n27, out3[5:0]}) );
  add_26_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_26_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in3[6:4], n23, in3[2], n22, in3[0]}), .SUM(out2) );
  add_26_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_26_DW01_add_4 add_30 ( .A({in2[6:4], n24, n25, in2[1:0]}), .B({in3[6:4], 
        n23, in3[2], n22, in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_26_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX2TH U1 ( .A(in3[1]), .Y(n22) );
  INVXLTH U2 ( .A(in2[4]), .Y(n19) );
  INVXLTH U4 ( .A(n19), .Y(n21) );
  CLKBUFX40 U3 ( .A(in3[3]), .Y(n23) );
  CLKBUFX40 U5 ( .A(in2[3]), .Y(n24) );
  CLKBUFX40 U6 ( .A(in2[2]), .Y(n25) );
  CLKBUFX40 U13 ( .A(n27), .Y(out3[6]) );
endmodule


module tc_sm_107 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U10 ( .A(in[5]), .Y(n27) );
  INVXLTH U11 ( .A(in[4]), .Y(n28) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_106 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n25, n26, n28, n29, n30, n31, n32,
         n33, n35;

  NAND3XL U3 ( .A(n28), .B(n29), .C(n6), .Y(out[1]) );
  OAI211XL U5 ( .A0(in[6]), .A1(n31), .B0(n5), .C0(n6), .Y(out[3]) );
  OR2X2 U6 ( .A(n30), .B(n8), .Y(n25) );
  OR2XLTH U7 ( .A(in[6]), .B(n32), .Y(n26) );
  NAND3XLTH U8 ( .A(n25), .B(n26), .C(n6), .Y(out[2]) );
  CLKINVX1 U9 ( .A(in[6]), .Y(n30) );
  OAI2B11X4 U10 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OAI21XL U11 ( .A0(n7), .A1(n31), .B0(in[6]), .Y(n5) );
  NOR3X1 U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  OR2X2 U13 ( .A(n30), .B(n10), .Y(n28) );
  AOI2BB1X4 U14 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n9) );
  INVXLTH U16 ( .A(in[3]), .Y(n31) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  OR2XLTH U18 ( .A(in[6]), .B(n33), .Y(n29) );
  XOR2XLTH U19 ( .A(in[0]), .B(n33), .Y(n10) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  INVXLTH U21 ( .A(in[2]), .Y(n32) );
  XOR2XLTH U22 ( .A(in[2]), .B(n9), .Y(n8) );
  INVXLTH U23 ( .A(in[1]), .Y(n33) );
  AO21X4 U4 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n35) );
  CLKINVX40 U24 ( .A(n35), .Y(n6) );
endmodule


module tc_sm_105 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n26, n27,
         n28;

  NAND2BXL U4 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211X2TH U5 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  CLKINVX1TH U6 ( .A(in[3]), .Y(n22) );
  OAI221X2TH U7 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2]) );
  OAI221X2TH U8 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1]) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U10 ( .A(in[6]), .Y(n19) );
  XNOR2XLTH U11 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U13 ( .A(in[2]), .Y(n23) );
  OAI21XLTH U14 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U16 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXL U19 ( .A(in[5]), .Y(n20) );
  INVXL U20 ( .A(in[4]), .Y(n21) );
  AOI33X4 U3 ( .A0(n21), .A1(n27), .A2(n20), .B0(n28), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U18 ( .A(n26), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n27) );
  AOI21BX4 U22 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n28) );
endmodule


module tc_sm_104 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n20, n21, n22, n23;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  CLKINVX1TH U3 ( .A(in[6]), .Y(n20) );
  OAI221XLTH U4 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n23), .C0(n6), .Y(out[1]) );
  OAI211XLTH U5 ( .A0(in[6]), .A1(n21), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI221XLTH U6 ( .A0(n20), .A1(n8), .B0(in[6]), .B1(n22), .C0(n6), .Y(out[2])
         );
  AOI21X8 U8 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n6) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  XOR2XLTH U10 ( .A(in[0]), .B(n23), .Y(n10) );
  INVXLTH U11 ( .A(in[1]), .Y(n23) );
  OAI21XLTH U12 ( .A0(n7), .A1(n21), .B0(in[6]), .Y(n5) );
  INVXLTH U13 ( .A(in[3]), .Y(n21) );
  INVXLTH U14 ( .A(in[2]), .Y(n22) );
  XOR2XLTH U15 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n9) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  AOI2BB1X2 U19 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
endmodule


module total_3_test_21 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n5, n6, n7, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_107 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_106 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_105 sm_tc_3 ( .out(c1), .in({c[4], n44, c[2:0]}) );
  sm_tc_104 sm_tc_4 ( .out(in1), .in(in) );
  add_26 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_107 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_106 tc_sm_2 ( .out(w6), .in({n5, w66[5:0]}) );
  tc_sm_105 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_104 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up2[1]) );
  SDFFRQX2TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n46), .CK(clk), .RN(n6), .Q(
        up1[0]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up3[0]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n53), .CK(clk), .RN(n7), .Q(
        h) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n54), .CK(clk), .RN(n6), 
        .Q(up2[0]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up2[2]) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up2[4]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n46), .CK(clk), .RN(n6), 
        .Q(up2[3]) );
  SDFFRQX4TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n50), .CK(clk), .RN(n7), 
        .Q(up1[4]) );
  SDFFRQX2TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up3[4]) );
  SDFFRQX4TH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n52), .CK(clk), .RN(n6), 
        .Q(up1[1]) );
  SDFFRQX2 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n53), .CK(clk), .RN(n6), 
        .Q(up1[2]) );
  BUFX10 U3 ( .A(w66[6]), .Y(n5) );
  CLKBUFX1TH U4 ( .A(rst), .Y(n7) );
  CLKBUFX4TH U5 ( .A(rst), .Y(n6) );
  SDFFRX4 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n54), .CK(clk), .RN(n6), 
        .Q(up3[2]) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up3[1]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n48), .CK(clk), .RN(n7), 
        .Q(up1[3]) );
  SDFFRX4 up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n52), .CK(clk), .RN(n6), 
        .Q(up3[3]) );
  CLKBUFX40 U38 ( .A(c[3]), .Y(n44) );
  DLY1X1TH U39 ( .A(n47), .Y(n45) );
  INVXLTH U40 ( .A(n47), .Y(n46) );
  DLY1X1TH U41 ( .A(n51), .Y(n47) );
  INVXLTH U42 ( .A(n47), .Y(n48) );
  INVXLTH U43 ( .A(n51), .Y(n49) );
  DLY1X1TH U44 ( .A(test_se), .Y(n50) );
  INVXLTH U45 ( .A(test_se), .Y(n51) );
  INVXLTH U46 ( .A(n45), .Y(n52) );
  INVXLTH U47 ( .A(n45), .Y(n53) );
  INVXLTH U48 ( .A(n47), .Y(n54) );
endmodule


module sm_tc_103 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n26, n27, n30;

  CLKBUFX2 U2 ( .A(in[4]), .Y(n22) );
  INVX4 U3 ( .A(n22), .Y(n26) );
  CLKBUFX1TH U5 ( .A(in[0]), .Y(out[0]) );
  OAI22XLTH U6 ( .A0(n22), .A1(n27), .B0(n5), .B1(n26), .Y(out[2]) );
  NOR2X4 U8 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI2BB2X4 U9 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n26), .Y(out[1]) );
  XNOR2X2 U10 ( .A(n27), .B(n8), .Y(n5) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  AOI31X2TH U12 ( .A0(n3), .A1(n4), .A2(n5), .B0(n26), .Y(out[4]) );
  XNOR2X4TH U13 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKINVX1TH U14 ( .A(in[2]), .Y(n27) );
  OAI2BB2XLTH U15 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[5]) );
  OAI2BB1X4 U4 ( .A0N(in[0]), .A1N(in[1]), .B0(n30), .Y(n6) );
  OR2X8 U7 ( .A(n30), .B(in[2]), .Y(n7) );
  CLKINVX40 U18 ( .A(n8), .Y(n30) );
endmodule


module sm_tc_102 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n4, n5, n6, n7, n8, n9, n24, n27, n28, n30, n31;

  OAI2BB2X1TH U3 ( .B0(n28), .B1(n7), .A0N(in[1]), .A1N(n28), .Y(out[1]) );
  OAI2BB2X1TH U4 ( .B0(n28), .B1(n5), .A0N(in[3]), .A1N(n28), .Y(out[3]) );
  AOI31X2TH U5 ( .A0(n4), .A1(n5), .A2(n6), .B0(n28), .Y(out[4]) );
  OAI22X2 U6 ( .A0(in[4]), .A1(n27), .B0(n28), .B1(n6), .Y(out[2]) );
  INVX6TH U7 ( .A(in[4]), .Y(n28) );
  CLKINVX1TH U8 ( .A(n24), .Y(out[6]) );
  XNOR2X1TH U10 ( .A(n8), .B(in[3]), .Y(n5) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n27) );
  INVXLTH U12 ( .A(out[4]), .Y(n24) );
  INVXLTH U13 ( .A(n24), .Y(out[5]) );
  NOR2BXLTH U14 ( .AN(n7), .B(in[0]), .Y(n4) );
  NAND2XLTH U15 ( .A(n9), .B(n27), .Y(n8) );
  BUFX2TH U16 ( .A(in[0]), .Y(out[0]) );
  XOR2X1 U2 ( .A(in[2]), .B(n9), .Y(n6) );
  AOI21BX4 U9 ( .A0(in[0]), .A1(in[1]), .B0N(n31), .Y(n30) );
  CLKINVX40 U17 ( .A(n30), .Y(n7) );
  OR2X8 U18 ( .A(in[1]), .B(in[0]), .Y(n31) );
  CLKINVX40 U19 ( .A(n31), .Y(n9) );
endmodule


module sm_tc_101 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n23, n24, n28, n29;

  AO21X2 U2 ( .A0(in[0]), .A1(n24), .B0(n8), .Y(n6) );
  NOR2X4 U3 ( .A(n24), .B(in[0]), .Y(n8) );
  BUFX6 U4 ( .A(in[4]), .Y(n23) );
  INVX2 U5 ( .A(n23), .Y(n28) );
  XNOR2X1TH U6 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX2 U7 ( .A(in[1]), .Y(n24) );
  AOI31X2TH U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n28), .Y(out[4]) );
  OAI2BB2X1 U9 ( .B0(n28), .B1(n6), .A0N(n24), .A1N(n28), .Y(out[1]) );
  CLKBUFX1TH U10 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X1TH U11 ( .B0(n28), .B1(n4), .A0N(in[3]), .A1N(n28), .Y(out[3]) );
  OAI22X4 U12 ( .A0(n23), .A1(n29), .B0(n28), .B1(n5), .Y(out[2]) );
  INVX2TH U13 ( .A(in[2]), .Y(n29) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  CLKNAND2X2TH U15 ( .A(n8), .B(n29), .Y(n7) );
  XNOR2X1TH U16 ( .A(n29), .B(n8), .Y(n5) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  BUFX2TH U18 ( .A(in[0]), .Y(out[0]) );
endmodule


module sm_tc_100 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  CLKINVX2TH U2 ( .A(out[4]), .Y(n18) );
  XNOR2X2TH U3 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX1TH U4 ( .A(n18), .Y(out[5]) );
  OAI2BB2X1TH U5 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U6 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U7 ( .A(n18), .Y(out[6]) );
  CLKINVX2TH U8 ( .A(in[4]), .Y(n22) );
  NOR2X3TH U9 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U10 ( .A(in[2]), .Y(n21) );
  AOI31X2TH U11 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U12 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI22X1TH U13 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  OAI2BB2X1TH U14 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  XNOR2X1TH U15 ( .A(n21), .B(n8), .Y(n5) );
  NAND2XLTH U16 ( .A(n8), .B(n21), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_25_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_25_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  NAND2X2 U1 ( .A(A[5]), .B(B[5]), .Y(n3) );
  NAND2X1 U3 ( .A(carry[5]), .B(B[5]), .Y(n4) );
  NAND3X4 U4 ( .A(n2), .B(n3), .C(n4), .Y(carry[6]) );
  CLKXOR2X1TH U6 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U7 ( .A(B[0]), .B(A[0]), .Y(n1) );
  AND2X8 U2 ( .A(A[5]), .B(carry[5]), .Y(n5) );
  CLKINVX40 U5 ( .A(n5), .Y(n2) );
  XNOR3X2 U8 ( .A(A[5]), .B(carry[5]), .C(B[5]), .Y(n6) );
  CLKINVX40 U9 ( .A(n6), .Y(SUM[5]) );
endmodule


module add_25_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR3X4TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_25_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX4TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X4 U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  XOR2XL U2 ( .A(A[6]), .B(B[6]), .Y(n2) );
  CLKXOR2X1TH U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_25_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2TH U1_3 ( .A(A[3]), .B(carry[3]), .CI(B[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3XL U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_25_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_25 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n19, n20, n21, n22, n23, n24, n25;

  add_25_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, n24, temp1_3_, temp1_2_, 
        temp1_1_, n25}), .B({in2[6:3], n23, in2[1:0]}), .SUM(out3) );
  add_25_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, n21, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_25_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, n24, temp1_3_, temp1_2_, 
        temp1_1_, n25}), .B({in3[6:2], n22, in3[0]}), .SUM(out2) );
  add_25_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, n24, temp1_3_, n20, 
        temp1_1_, n25}), .B({temp2_6_, temp2_5_, n21, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_25_DW01_add_4 add_30 ( .A({in2[6:3], n23, in2[1:0]}), .B({in3[6:2], n22, 
        in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_25_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX1 U1 ( .A(in3[1]), .Y(n22) );
  CLKBUFX2 U2 ( .A(temp2_4_), .Y(n21) );
  CLKBUFX1TH U3 ( .A(in2[2]), .Y(n23) );
  INVXLTH U4 ( .A(temp1_2_), .Y(n19) );
  INVXLTH U5 ( .A(n19), .Y(n20) );
  CLKBUFX40 U6 ( .A(temp1_4_), .Y(n24) );
  CLKBUFX40 U13 ( .A(temp1_0_), .Y(n25) );
endmodule


module tc_sm_103 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n28) );
  XNOR2XLTH U7 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(in[6]), .Y(n24) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n26) );
  INVXLTH U12 ( .A(in[5]), .Y(n25) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n27) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U16 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_102 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n7, n8, n9, n10, n11, n12, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n35, n36, n37, n38, n40;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[5]), .C0(in[4]), .Y(n11) );
  NAND2XL U3 ( .A(n33), .B(n29), .Y(out[3]) );
  NOR2X2 U4 ( .A(n35), .B(n10), .Y(n24) );
  NOR2XLTH U5 ( .A(in[6]), .B(n38), .Y(n25) );
  INVXLTH U6 ( .A(n29), .Y(n26) );
  OR3X2 U8 ( .A(n24), .B(n25), .C(n26), .Y(out[1]) );
  AOI21X8 U9 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n29) );
  NAND2X2 U10 ( .A(n29), .B(n31), .Y(n27) );
  NAND2X3 U11 ( .A(n30), .B(n28), .Y(out[2]) );
  CLKINVX4 U12 ( .A(n27), .Y(n28) );
  INVXLTH U13 ( .A(in[6]), .Y(n35) );
  OR2X2 U14 ( .A(n35), .B(n8), .Y(n30) );
  OR2XLTH U15 ( .A(in[6]), .B(n37), .Y(n31) );
  OR2X1TH U16 ( .A(n7), .B(n36), .Y(n32) );
  OA21X1 U18 ( .A0(in[6]), .A1(n36), .B0(n5), .Y(n33) );
  INVXLTH U19 ( .A(in[3]), .Y(n36) );
  AOI2BB1X4 U20 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  NOR3X1TH U21 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  XOR2XLTH U22 ( .A(in[0]), .B(n38), .Y(n10) );
  INVXLTH U23 ( .A(in[1]), .Y(n38) );
  NAND2BXLTH U24 ( .AN(in[0]), .B(n29), .Y(out[0]) );
  INVXLTH U25 ( .A(in[2]), .Y(n37) );
  XOR2XLTH U26 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U27 ( .A(in[0]), .B(in[1]), .Y(n9) );
  CLKBUFX1TH U28 ( .A(in[6]), .Y(out[4]) );
  AND2X8 U17 ( .A(n32), .B(in[6]), .Y(n40) );
  CLKINVX40 U29 ( .A(n40), .Y(n5) );
endmodule


module tc_sm_101 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n23, n24, n25, n27, n28, n29,
         n30, n31, n32, n33;

  OAI221X1TH U3 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[2]) );
  OAI221XL U4 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[1])
         );
  OAI211XLTH U5 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
  INVX2TH U7 ( .A(in[5]), .Y(n21) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n23) );
  INVXLTH U9 ( .A(in[6]), .Y(n20) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U13 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U15 ( .A(in[2]), .Y(n24) );
  OAI21XLTH U16 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  INVXLTH U17 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  DLY1X1TH U6 ( .A(in[4]), .Y(n27) );
  AOI33X4 U10 ( .A0(n29), .A1(n30), .A2(n31), .B0(n33), .B1(n32), .B2(in[4]), 
        .Y(n28) );
  CLKINVX40 U20 ( .A(n28), .Y(n8) );
  CLKINVX40 U21 ( .A(n27), .Y(n29) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n30) );
  CLKINVX40 U23 ( .A(in[5]), .Y(n31) );
  CLKINVX40 U24 ( .A(n21), .Y(n32) );
  AOI21BX4 U25 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n33) );
endmodule


module tc_sm_100 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n19, n21, n22, n23, n24, n25, n26;

  OAI221XL U3 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n25), .C0(n19), .Y(out[2])
         );
  OAI211XLTH U4 ( .A0(in[6]), .A1(n24), .B0(n7), .C0(n19), .Y(out[3]) );
  INVXLTH U5 ( .A(in[6]), .Y(n21) );
  BUFX5 U6 ( .A(n8), .Y(n19) );
  INVX1TH U7 ( .A(in[3]), .Y(n24) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  NAND2BXLTH U9 ( .AN(in[0]), .B(n19), .Y(out[0]) );
  OAI221XLTH U10 ( .A0(n21), .A1(n12), .B0(in[6]), .B1(n26), .C0(n19), .Y(
        out[1]) );
  CLKBUFX1TH U11 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U12 ( .A0(n9), .A1(n24), .B0(in[6]), .Y(n7) );
  XNOR2XLTH U13 ( .A(n25), .B(n11), .Y(n10) );
  INVXLTH U14 ( .A(in[2]), .Y(n25) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI2BB1X4 U18 ( .A0N(n24), .A1N(n9), .B0(in[6]), .Y(n13) );
  INVX2 U19 ( .A(in[5]), .Y(n22) );
  OAI33X4 U20 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n22), .B2(
        n23), .Y(n8) );
  INVXL U21 ( .A(in[4]), .Y(n23) );
endmodule


module total_3_test_22 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n64, w5_4_, n7, n8, n9, n10, n45, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_103 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_102 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_101 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_100 sm_tc_4 ( .out(in1), .in(in) );
  add_25 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_103 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_102 tc_sm_2 ( .out(w6), .in({n8, w66[5:0]}) );
  tc_sm_101 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_100 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n50), .CK(clk), .RN(n9), 
        .Q(up1[4]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n57), .CK(clk), .RN(n10), 
        .Q(h) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n49), .CK(clk), .RN(n9), 
        .Q(up3[2]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n54), .CK(clk), .RN(n9), 
        .Q(n64) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n54), .CK(clk), .RN(n9), 
        .Q(up2[1]) );
  SDFFRQX2TH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n49), .CK(clk), .RN(n9), 
        .Q(up2[2]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n58), .CK(clk), .RN(n9), 
        .Q(up2[0]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n53), .CK(clk), .RN(n10), 
        .Q(up1[3]) );
  SDFFRQX2 up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n57), .CK(clk), .RN(n9), 
        .Q(up3[4]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n50), .CK(clk), .RN(n9), 
        .Q(up3[0]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n59), .CK(clk), .RN(n9), 
        .Q(up1[2]) );
  SDFFRQX2 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n56), .CK(clk), .RN(n9), 
        .Q(up1[1]) );
  SDFFRQX2 up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n58), .CK(clk), .RN(n10), 
        .Q(up2[4]) );
  INVX20 U3 ( .A(n7), .Y(n8) );
  CLKINVX12 U4 ( .A(w66[6]), .Y(n7) );
  CLKBUFX1TH U5 ( .A(rst), .Y(n10) );
  CLKBUFX4TH U6 ( .A(rst), .Y(n9) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n53), .CK(clk), .RN(n9), 
        .Q(up3[1]) );
  SDFFRX4 up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n59), .CK(clk), .RN(n9), .Q(
        up1[0]) );
  SDFFRX4 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n56), .CK(clk), .RN(n9), 
        .Q(n45) );
  INVXLTH U39 ( .A(n52), .Y(n49) );
  INVXLTH U40 ( .A(n51), .Y(n50) );
  DLY1X1TH U41 ( .A(n55), .Y(n51) );
  DLY1X1TH U42 ( .A(n55), .Y(n52) );
  INVXLTH U43 ( .A(n52), .Y(n53) );
  INVXLTH U44 ( .A(n51), .Y(n54) );
  INVXLTH U45 ( .A(test_se), .Y(n55) );
  INVXLTH U46 ( .A(n52), .Y(n56) );
  INVXLTH U47 ( .A(n51), .Y(n57) );
  INVXLTH U48 ( .A(n52), .Y(n58) );
  INVXLTH U49 ( .A(n51), .Y(n59) );
  DLY1X1TH U50 ( .A(n45), .Y(up2[3]) );
  DLY1X1TH U51 ( .A(n64), .Y(up3[3]) );
endmodule


module sm_tc_99 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n23, n26, n27;

  AO21X1 U2 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  DLY2X1TH U3 ( .A(in[0]), .Y(out[0]) );
  XNOR2X4TH U4 ( .A(n23), .B(n8), .Y(n5) );
  CLKBUFX1TH U6 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X1TH U7 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  AOI31X2TH U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  OAI22X1TH U9 ( .A0(in[4]), .A1(n23), .B0(n22), .B1(n5), .Y(out[2]) );
  XNOR2X2TH U10 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX6TH U11 ( .A(in[4]), .Y(n22) );
  OAI2BB2X2TH U12 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKINVX1TH U14 ( .A(in[2]), .Y(n23) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  AND2X8 U5 ( .A(n8), .B(n23), .Y(n26) );
  CLKINVX40 U13 ( .A(n26), .Y(n7) );
  OR2X8 U17 ( .A(in[1]), .B(in[0]), .Y(n27) );
  CLKINVX40 U18 ( .A(n27), .Y(n8) );
endmodule


module sm_tc_98 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n28, n31, n32;

  NAND2X2 U2 ( .A(n21), .B(n22), .Y(n24) );
  NAND2X2 U3 ( .A(n8), .B(n31), .Y(n7) );
  OAI2BB2X1 U4 ( .B0(n32), .B1(n4), .A0N(in[3]), .A1N(n32), .Y(out[3]) );
  INVX2 U5 ( .A(n26), .Y(n32) );
  NOR2X4 U6 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKNAND2X2 U7 ( .A(n23), .B(n24), .Y(n4) );
  NAND3XLTH U8 ( .A(n3), .B(n4), .C(n5), .Y(n25) );
  OAI2BB2X2 U9 ( .B0(n32), .B1(n6), .A0N(in[1]), .A1N(n32), .Y(out[1]) );
  INVX2 U10 ( .A(n28), .Y(out[5]) );
  BUFX6 U11 ( .A(in[4]), .Y(n26) );
  AO21XL U12 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  INVXLTH U13 ( .A(n7), .Y(n21) );
  CLKNAND2X2TH U14 ( .A(n19), .B(n20), .Y(n5) );
  NAND2XLTH U15 ( .A(n17), .B(n18), .Y(n20) );
  NAND2XLTH U16 ( .A(n31), .B(n8), .Y(n19) );
  CLKINVX1TH U17 ( .A(n31), .Y(n17) );
  INVXLTH U18 ( .A(n8), .Y(n18) );
  INVX2TH U19 ( .A(in[2]), .Y(n31) );
  OAI22X4 U20 ( .A0(n26), .A1(n31), .B0(n32), .B1(n5), .Y(out[2]) );
  NAND2X2 U21 ( .A(n7), .B(in[3]), .Y(n23) );
  INVXLTH U22 ( .A(in[3]), .Y(n22) );
  AND2X2 U23 ( .A(n25), .B(n26), .Y(out[4]) );
  INVXLTH U24 ( .A(out[4]), .Y(n28) );
  NOR2BXLTH U25 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U26 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U27 ( .A(n28), .Y(out[6]) );
endmodule


module sm_tc_97 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n4, n5, n6, n7, n8, n9, n31, n32;

  DLY1X1TH U2 ( .A(in[0]), .Y(out[0]) );
  XNOR2X4 U3 ( .A(n31), .B(n9), .Y(n6) );
  INVX3TH U4 ( .A(in[4]), .Y(n32) );
  OAI22X2 U5 ( .A0(in[4]), .A1(n31), .B0(n32), .B1(n6), .Y(out[2]) );
  OAI2BB2X2 U6 ( .B0(n32), .B1(n7), .A0N(in[1]), .A1N(n32), .Y(out[1]) );
  AOI31X2 U7 ( .A0(n4), .A1(n5), .A2(n6), .B0(n32), .Y(out[4]) );
  OAI2BB2X2TH U8 ( .B0(n32), .B1(n5), .A0N(in[3]), .A1N(n32), .Y(out[3]) );
  XNOR2X1TH U9 ( .A(n8), .B(in[3]), .Y(n5) );
  CLKBUFX1TH U10 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  CLKINVX1TH U12 ( .A(in[2]), .Y(n31) );
  AO21X2 U13 ( .A0(in[0]), .A1(in[1]), .B0(n9), .Y(n7) );
  NOR2X4 U14 ( .A(in[1]), .B(in[0]), .Y(n9) );
  NAND2XLTH U15 ( .A(n9), .B(n31), .Y(n8) );
  NOR2BXLTH U16 ( .AN(n7), .B(in[0]), .Y(n4) );
endmodule


module sm_tc_96 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  CLKNAND2X2TH U2 ( .A(n8), .B(n21), .Y(n7) );
  OAI22X2TH U3 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  CLKINVX2 U4 ( .A(out[4]), .Y(n18) );
  XNOR2X1TH U5 ( .A(n21), .B(n8), .Y(n5) );
  NOR2X1TH U6 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U7 ( .A(in[2]), .Y(n21) );
  XNOR2X1TH U8 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKINVX2TH U9 ( .A(in[4]), .Y(n22) );
  AOI31X2TH U10 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U11 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U12 ( .A(n18), .Y(out[5]) );
  INVXLTH U13 ( .A(n18), .Y(out[6]) );
  CLKBUFX1TH U14 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X2TH U15 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  OAI2BB2XL U16 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_24_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X8 U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  CLKXOR2X2TH U2 ( .A(B[6]), .B(A[6]), .Y(n2) );
  CLKXOR2X1TH U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_24_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [6:2] carry;

  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKNAND2X2 U1 ( .A(n2), .B(n7), .Y(n8) );
  NAND2X1 U2 ( .A(n6), .B(carry[3]), .Y(n9) );
  NAND2X2 U3 ( .A(n8), .B(n9), .Y(SUM[3]) );
  CLKINVX2 U4 ( .A(n2), .Y(n6) );
  INVXLTH U5 ( .A(carry[3]), .Y(n7) );
  NAND2XL U6 ( .A(carry[3]), .B(B[3]), .Y(n4) );
  XOR2X1TH U7 ( .A(B[3]), .B(A[3]), .Y(n2) );
  NAND2XLTH U8 ( .A(A[3]), .B(B[3]), .Y(n5) );
  NAND2XLTH U9 ( .A(carry[3]), .B(A[3]), .Y(n3) );
  CLKAND2X2 U10 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U11 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND3X2TH U12 ( .A(n3), .B(n4), .C(n5), .Y(carry[4]) );
  XNOR3X2 U13 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n10) );
  CLKINVX40 U14 ( .A(n10), .Y(SUM[6]) );
endmodule


module add_24_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX2TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X8 U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  XOR2X1TH U2 ( .A(B[6]), .B(A[6]), .Y(n2) );
  CLKXOR2X1TH U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_24_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n3;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n3) );
endmodule


module add_24_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7;
  wire   [6:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n5), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  NAND2X2 U1 ( .A(n4), .B(n3), .Y(n6) );
  CLKNAND2X4 U2 ( .A(n2), .B(n7), .Y(carry[3]) );
  INVX3 U3 ( .A(n6), .Y(n7) );
  NAND2X2 U4 ( .A(carry[2]), .B(B[2]), .Y(n2) );
  XOR2X2 U5 ( .A(A[2]), .B(B[2]), .Y(n1) );
  CLKNAND2X2 U6 ( .A(carry[2]), .B(A[2]), .Y(n3) );
  AND2XLTH U7 ( .A(B[0]), .B(A[0]), .Y(n5) );
  CLKXOR2X1TH U8 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X2TH U9 ( .A(n1), .B(carry[2]), .Y(SUM[2]) );
  NAND2XLTH U10 ( .A(B[2]), .B(A[2]), .Y(n4) );
endmodule


module add_24_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n4, n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR2X3TH U1 ( .A(B[0]), .B(A[0]), .Y(n4) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKINVX40 U3 ( .A(n4), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[0]) );
endmodule


module add_24 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n21, n22, n23, n24, n25, n26, n27;

  add_24_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n27, temp1_0_}), .B(in2), .SUM(out3) );
  add_24_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, n26, 
        temp2_1_, temp2_0_}), .B({in[6:3], n23, in[1:0]}), .SUM(out1) );
  add_24_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in3[6:3], n25, n24, n22}), .SUM(
        out2) );
  add_24_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n21, 
        n27, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, n26, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_24_DW01_add_4 add_30 ( .A(in2), .B({in3[6:3], n25, in3[1], n22}), .SUM({
        temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_})
         );
  add_24_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX2TH U1 ( .A(temp1_2_), .Y(n21) );
  BUFX10 U2 ( .A(in3[0]), .Y(n22) );
  CLKBUFX1TH U3 ( .A(in3[1]), .Y(n24) );
  CLKBUFX1TH U4 ( .A(in[2]), .Y(n23) );
  BUFX2TH U5 ( .A(in3[2]), .Y(n25) );
  BUFX8 U6 ( .A(temp2_2_), .Y(n26) );
  CLKBUFX40 U13 ( .A(temp1_1_), .Y(n27) );
endmodule


module tc_sm_99 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n25, n27, n28, n29, n30, n31, n32;

  CLKBUFX2TH U3 ( .A(in[6]), .Y(n25) );
  INVXLTH U4 ( .A(in[1]), .Y(n32) );
  INVXLTH U5 ( .A(in[2]), .Y(n31) );
  XNOR2XLTH U6 ( .A(n31), .B(n11), .Y(n10) );
  OAI33X4TH U7 ( .A0(in[4]), .A1(n25), .A2(in[5]), .B0(n13), .B1(n28), .B2(n29), .Y(n8) );
  INVXLTH U8 ( .A(in[4]), .Y(n29) );
  INVXLTH U9 ( .A(in[5]), .Y(n28) );
  CLKINVX1TH U10 ( .A(in[3]), .Y(n30) );
  CLKBUFX1TH U11 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U12 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(n25), .Y(n27) );
  OAI221XLTH U17 ( .A0(n27), .A1(n12), .B0(n25), .B1(n32), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U18 ( .A0(n27), .A1(n10), .B0(n25), .B1(n31), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U19 ( .A0(n9), .A1(n30), .B0(n25), .Y(n7) );
  OAI211XLTH U20 ( .A0(n25), .A1(n30), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U21 ( .A0N(n30), .A1N(n9), .B0(n25), .Y(n13) );
endmodule


module tc_sm_98 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n25, n26, n27, n28, n29, n30, n32,
         n33, n34, n35, n36, n37, n39;

  INVX2 U3 ( .A(in[3]), .Y(n35) );
  OAI33X4 U5 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n34), .B2(n33), .Y(n8) );
  OAI2BB1X2 U6 ( .A0N(n35), .A1N(n9), .B0(in[6]), .Y(n13) );
  NAND3X1 U7 ( .A(n25), .B(n26), .C(n30), .Y(out[2]) );
  INVX2TH U8 ( .A(in[4]), .Y(n34) );
  OAI21X3TH U9 ( .A0(n9), .A1(n35), .B0(in[6]), .Y(n7) );
  OR2X1 U10 ( .A(n32), .B(n10), .Y(n25) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  OR2XLTH U12 ( .A(in[6]), .B(n36), .Y(n26) );
  NAND2XLTH U13 ( .A(n29), .B(n30), .Y(out[3]) );
  OA21XLTH U14 ( .A0(in[6]), .A1(n35), .B0(n7), .Y(n29) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n30), .Y(out[0]) );
  OR2XLTH U16 ( .A(n32), .B(n12), .Y(n27) );
  OR2XLTH U17 ( .A(in[6]), .B(n37), .Y(n28) );
  CLKBUFX1TH U18 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U19 ( .A(n36), .B(n11), .Y(n10) );
  BUFX10 U20 ( .A(n8), .Y(n30) );
  INVX2 U21 ( .A(in[5]), .Y(n33) );
  INVXLTH U22 ( .A(in[1]), .Y(n37) );
  XNOR2XLTH U23 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U24 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U25 ( .A(in[2]), .Y(n36) );
  INVXL U26 ( .A(in[6]), .Y(n32) );
  AND3X8 U4 ( .A(n27), .B(n28), .C(n30), .Y(n39) );
  CLKINVX40 U27 ( .A(n39), .Y(out[1]) );
endmodule


module tc_sm_97 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n19, n20, n21, n22, n23, n24, n26,
         n27;

  OAI211X1 U3 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n27), .Y(out[3]) );
  NAND2BXL U4 ( .AN(in[0]), .B(n27), .Y(out[0]) );
  OAI221X2TH U5 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n27), .Y(
        out[1]) );
  OAI221X2TH U6 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n27), .Y(
        out[2]) );
  INVXLTH U7 ( .A(in[6]), .Y(n19) );
  CLKBUFX1TH U8 ( .A(in[6]), .Y(out[4]) );
  OAI33X4 U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n20), .B2(n21), .Y(n8) );
  OAI2BB1X4 U10 ( .A0N(n22), .A1N(n9), .B0(in[6]), .Y(n13) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n22) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U13 ( .A(in[4]), .Y(n21) );
  INVXLTH U14 ( .A(in[5]), .Y(n20) );
  INVXLTH U15 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U17 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U19 ( .A(in[2]), .Y(n23) );
  OAI21XLTH U20 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  CLKINVX40 U21 ( .A(n8), .Y(n26) );
  CLKINVX40 U22 ( .A(n26), .Y(n27) );
endmodule


module tc_sm_96 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n23, n24, n25, n27, n28, n29,
         n30, n31;

  OAI221X2TH U3 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[2]) );
  OAI221X1 U4 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[1])
         );
  OAI211XL U5 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
  CLKBUFX1TH U6 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U9 ( .A(in[6]), .Y(n20) );
  CLKINVX1TH U10 ( .A(in[3]), .Y(n23) );
  INVXLTH U12 ( .A(in[5]), .Y(n21) );
  XNOR2XLTH U13 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U15 ( .A(in[2]), .Y(n24) );
  INVXLTH U16 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI21XLTH U19 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  NOR3X1TH U20 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U7 ( .A(n29), .Y(n27) );
  AOI33X4 U8 ( .A0(n29), .A1(n30), .A2(n21), .B0(n31), .B1(in[5]), .B2(n27), 
        .Y(n28) );
  CLKINVX40 U11 ( .A(n28), .Y(n8) );
  CLKINVX40 U21 ( .A(in[4]), .Y(n29) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n30) );
  AOI21BX4 U23 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n31) );
endmodule


module total_3_test_23 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n4, n5, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_99 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_98 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_97 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_96 sm_tc_4 ( .out(in1), .in(in) );
  add_24 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_99 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_98 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_97 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_96 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up3[3]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n43), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n46), .CK(clk), .RN(n5), .Q(
        h) );
  SDFFRQXLTH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n43), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n46), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n45), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  SDFFRQX1TH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up1[2]) );
  SDFFRQXLTH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n47), .CK(clk), .RN(n5), .Q(
        up1[0]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRQXL up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n45), .CK(clk), .RN(n4), 
        .Q(up1[1]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRQX2 up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n5) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n4) );
  SDFFRX4 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up2[3]) );
  DLY1X1TH U37 ( .A(n44), .Y(n42) );
  INVXLTH U38 ( .A(n44), .Y(n43) );
  DLY1X1TH U39 ( .A(n48), .Y(n44) );
  INVXLTH U40 ( .A(n44), .Y(n45) );
  INVXLTH U41 ( .A(n48), .Y(n46) );
  DLY1X1TH U42 ( .A(test_se), .Y(n47) );
  INVXLTH U43 ( .A(test_se), .Y(n48) );
  INVXLTH U44 ( .A(n42), .Y(n49) );
  INVXLTH U45 ( .A(n42), .Y(n50) );
  INVXLTH U46 ( .A(n44), .Y(n51) );
endmodule


module sm_tc_95 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n19, n20, n24, n25, n28, n29, n30, n31;

  AOI31X2 U3 ( .A0(n3), .A1(n28), .A2(n5), .B0(n25), .Y(out[4]) );
  XNOR2X2 U4 ( .A(n24), .B(n8), .Y(n5) );
  BUFX8 U5 ( .A(in[1]), .Y(n19) );
  BUFX8 U7 ( .A(in[4]), .Y(n20) );
  INVX2 U8 ( .A(in[2]), .Y(n24) );
  AO21X2 U10 ( .A0(n31), .A1(n19), .B0(n8), .Y(n6) );
  NOR2X4 U11 ( .A(n19), .B(n31), .Y(n8) );
  INVX10 U12 ( .A(n20), .Y(n25) );
  OAI2BB2X1TH U13 ( .B0(n25), .B1(n28), .A0N(in[3]), .A1N(n25), .Y(out[3]) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX2TH U15 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U18 ( .AN(n6), .B(n31), .Y(n3) );
  CLKBUFX40 U2 ( .A(n4), .Y(n28) );
  AO2B2BX4 U6 ( .A0(n25), .A1N(n24), .B0(n29), .B1N(n25), .Y(out[2]) );
  CLKINVX40 U9 ( .A(n5), .Y(n29) );
  AO2B2X4 U16 ( .B0(n19), .B1(n25), .A0(n20), .A1N(n6), .Y(out[1]) );
  AND2X8 U19 ( .A(n24), .B(n8), .Y(n30) );
  XOR2X1 U20 ( .A(n30), .B(in[3]), .Y(n4) );
  CLKBUFX40 U21 ( .A(in[0]), .Y(n31) );
endmodule


module sm_tc_94 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n19, n20, n21, n22, n23, n24, n26, n29,
         n30, n33, n34;

  INVX4 U3 ( .A(in[4]), .Y(n29) );
  CLKNAND2X2TH U4 ( .A(n7), .B(in[3]), .Y(n23) );
  INVX2TH U5 ( .A(in[2]), .Y(n30) );
  OAI2BB2X4 U6 ( .B0(n29), .B1(n6), .A0N(in[1]), .A1N(n29), .Y(out[1]) );
  INVX2 U7 ( .A(n7), .Y(n21) );
  AOI31X4TH U9 ( .A0(n3), .A1(n4), .A2(n5), .B0(n29), .Y(out[4]) );
  OAI2BB2X1TH U10 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  NAND2X3 U11 ( .A(n30), .B(n8), .Y(n19) );
  NAND2X5 U12 ( .A(n17), .B(n34), .Y(n20) );
  CLKNAND2X12 U13 ( .A(n19), .B(n20), .Y(n5) );
  CLKINVX2TH U14 ( .A(n30), .Y(n17) );
  CLKNAND2X4 U16 ( .A(n21), .B(n22), .Y(n24) );
  NAND2X8 U17 ( .A(n23), .B(n24), .Y(n4) );
  INVX3TH U18 ( .A(in[3]), .Y(n22) );
  INVXLTH U19 ( .A(out[4]), .Y(n26) );
  INVXLTH U20 ( .A(n26), .Y(out[5]) );
  INVXLTH U21 ( .A(n26), .Y(out[6]) );
  AO21X2 U22 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2BXLTH U23 ( .AN(n6), .B(in[0]), .Y(n3) );
  BUFX2TH U25 ( .A(in[0]), .Y(out[0]) );
  NAND2BX8 U2 ( .AN(n34), .B(n30), .Y(n7) );
  AO2B2BX4 U8 ( .A0(n29), .A1N(n30), .B0(n33), .B1N(n5), .Y(out[2]) );
  CLKINVX40 U15 ( .A(n29), .Y(n33) );
  OR2X8 U24 ( .A(in[1]), .B(in[0]), .Y(n34) );
  CLKINVX40 U26 ( .A(n34), .Y(n8) );
endmodule


module sm_tc_93 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n20, n21, n24;

  OAI22X4 U2 ( .A0(in[4]), .A1(n20), .B0(n21), .B1(n5), .Y(out[2]) );
  XNOR2X1 U3 ( .A(n20), .B(n8), .Y(n5) );
  AOI31X2 U5 ( .A0(n3), .A1(n4), .A2(n5), .B0(n21), .Y(out[4]) );
  XNOR2X1 U6 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX2 U7 ( .A(in[4]), .Y(n21) );
  OAI2BB2X1 U8 ( .B0(n21), .B1(n4), .A0N(in[3]), .A1N(n21), .Y(out[3]) );
  NAND2XLTH U9 ( .A(n8), .B(n20), .Y(n7) );
  NOR2X2TH U10 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n20) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U13 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[6]) );
  AO21X2 U15 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  AO2B2X4 U4 ( .B0(in[1]), .B1(n21), .A0(n24), .A1N(n21), .Y(out[1]) );
  CLKINVX40 U17 ( .A(n6), .Y(n24) );
endmodule


module sm_tc_92 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  OAI2BB2X2 U5 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  AO21X2 U2 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2BX1 U3 ( .AN(n6), .B(in[0]), .Y(n3) );
  AOI31X1 U4 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NAND2X2 U6 ( .A(n8), .B(n21), .Y(n7) );
  INVX1TH U7 ( .A(out[4]), .Y(n18) );
  CLKBUFX1TH U8 ( .A(in[0]), .Y(out[0]) );
  NOR2X2TH U9 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X1TH U10 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI22X1TH U11 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  INVXLTH U12 ( .A(n18), .Y(out[6]) );
  OAI2BB2X1TH U13 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  CLKINVX2TH U14 ( .A(in[4]), .Y(n22) );
  CLKINVX1TH U15 ( .A(in[2]), .Y(n21) );
  INVXLTH U16 ( .A(n18), .Y(out[5]) );
  XNOR2X1TH U17 ( .A(n21), .B(n8), .Y(n5) );
endmodule


module add_23_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X8TH U2 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  XOR2X3 U3 ( .A(B[6]), .B(A[6]), .Y(n2) );
  CLKAND2X2 U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_23_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_23_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_23_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n6, n1, n3, n4;
  wire   [6:2] carry;

  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR2X4TH U2 ( .A(n3), .B(carry[6]), .Y(n6) );
  XNOR2XLTH U3 ( .A(A[6]), .B(B[6]), .Y(n3) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKINVX40 U5 ( .A(n6), .Y(n4) );
  CLKINVX40 U6 ( .A(n4), .Y(SUM[6]) );
endmodule


module add_23_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(n1), .B(A[1]), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX1TH U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_23_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [6:2] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X2 U2 ( .A(B[1]), .B(n1), .C(A[1]), .Y(SUM[1]) );
  CLKNAND2X2 U3 ( .A(B[1]), .B(n1), .Y(n2) );
  CLKNAND2X2 U4 ( .A(B[1]), .B(A[1]), .Y(n3) );
  CLKNAND2X2 U5 ( .A(n1), .B(A[1]), .Y(n4) );
  CLKXOR2X2TH U7 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X8 U1 ( .A(B[0]), .B(A[0]), .Y(n5) );
  CLKINVX40 U6 ( .A(n5), .Y(n1) );
  AND3X8 U8 ( .A(n2), .B(n3), .C(n4), .Y(n6) );
  CLKINVX40 U9 ( .A(n6), .Y(carry[2]) );
endmodule


module add_23 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n21, n22, n23, n24;

  add_23_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n22, n23, 
        temp1_1_, n24}), .B(in2), .SUM(out3) );
  add_23_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_23_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n22, n23, 
        temp1_1_, n24}), .B(in3), .SUM(out2) );
  add_23_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n22, n23, 
        temp1_1_, n24}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, n21, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_23_DW01_add_4 add_30 ( .A(in2), .B(in3), .SUM({temp2_6_, temp2_5_, 
        temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_23_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2TH U1 ( .A(temp2_2_), .Y(n21) );
  CLKBUFX40 U2 ( .A(temp1_3_), .Y(n22) );
  CLKBUFX40 U3 ( .A(temp1_2_), .Y(n23) );
  CLKBUFX40 U4 ( .A(temp1_0_), .Y(n24) );
endmodule


module tc_sm_95 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n28) );
  XNOR2XLTH U7 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXLTH U10 ( .A(in[5]), .Y(n25) );
  INVXLTH U11 ( .A(in[4]), .Y(n26) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n27) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n24) );
  OAI21XLTH U16 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  OAI221XLTH U17 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U18 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(
        out[2]) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_94 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n20, n21, n23, n24, n25, n26;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OAI211XL U3 ( .A0(in[6]), .A1(n24), .B0(n5), .C0(n21), .Y(out[3]) );
  INVX12 U4 ( .A(n20), .Y(n21) );
  OAI221X1 U5 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n26), .C0(n21), .Y(out[1])
         );
  OAI221XL U6 ( .A0(n23), .A1(n8), .B0(in[6]), .B1(n25), .C0(n21), .Y(out[2])
         );
  AOI2BB1X4 U8 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  INVXLTH U9 ( .A(in[6]), .Y(n23) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  INVXLTH U11 ( .A(in[2]), .Y(n25) );
  XOR2XLTH U12 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n9) );
  XOR2XLTH U14 ( .A(in[0]), .B(n26), .Y(n10) );
  INVXLTH U15 ( .A(in[1]), .Y(n26) );
  OAI21XLTH U16 ( .A0(n7), .A1(n24), .B0(in[6]), .Y(n5) );
  INVXLTH U17 ( .A(in[3]), .Y(n24) );
  CLKBUFX1TH U18 ( .A(in[6]), .Y(out[4]) );
  INVX4 U19 ( .A(n6), .Y(n20) );
  AOI21X1 U20 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n6) );
  NAND2BXLTH U21 ( .AN(in[0]), .B(n21), .Y(out[0]) );
endmodule


module tc_sm_93 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n19, n20, n21, n22, n24, n25,
         n26, n27, n28, n29;

  OAI211XL U3 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n22), .Y(out[3]) );
  OR2X2 U4 ( .A(n24), .B(n10), .Y(n18) );
  OR2XLTH U5 ( .A(in[6]), .B(n28), .Y(n19) );
  NAND3XL U6 ( .A(n18), .B(n19), .C(n22), .Y(out[2]) );
  OR2X2 U7 ( .A(n24), .B(n12), .Y(n20) );
  OR2XLTH U8 ( .A(in[6]), .B(n29), .Y(n21) );
  NAND3XL U9 ( .A(n20), .B(n21), .C(n22), .Y(out[1]) );
  OAI2BB1X1 U10 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
  BUFX10 U11 ( .A(n8), .Y(n22) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n27) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U14 ( .A(in[6]), .Y(n24) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U16 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  XNOR2XLTH U17 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U19 ( .A(in[2]), .Y(n28) );
  INVXLTH U20 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U22 ( .AN(in[0]), .B(n22), .Y(out[0]) );
  OAI33X4 U23 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXL U24 ( .A(in[5]), .Y(n25) );
  INVXL U25 ( .A(in[4]), .Y(n26) );
endmodule


module tc_sm_92 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n20, n21, n22, n23, n24, n25,
         n27;

  OAI211XL U3 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n18), .Y(out[3]) );
  BUFX8 U4 ( .A(n8), .Y(n18) );
  OAI221XL U5 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n18), .Y(out[2])
         );
  OAI221XL U7 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n18), .Y(out[1])
         );
  INVXLTH U8 ( .A(in[6]), .Y(n20) );
  CLKBUFX1TH U9 ( .A(in[6]), .Y(out[4]) );
  CLKINVX1TH U10 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U12 ( .A(in[4]), .Y(n22) );
  XNOR2XLTH U13 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U15 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U17 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  INVX2 U18 ( .A(in[5]), .Y(n21) );
  INVXLTH U19 ( .A(in[2]), .Y(n24) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  OAI33X4 U21 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n21), .B2(
        n22), .Y(n8) );
  AO21X4 U6 ( .A0(n23), .A1(n9), .B0(n27), .Y(n13) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n27) );
endmodule


module total_3_test_24 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n66, n67, w5_4_, n4, n5, n6, n44, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_95 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_94 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_93 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_92 sm_tc_4 ( .out(in1), .in(in) );
  add_23 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2({b1[6:2], n4, b1[0]}), .in3(c1), .in(in1) );
  tc_sm_95 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_94 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_93 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_92 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up1[3]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n54), .CK(clk), .RN(n5), 
        .Q(n67) );
  SDFFRQX1TH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up1[1]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n52), .CK(clk), .RN(n6), .Q(
        h) );
  SDFFRQXLTH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n50), .CK(clk), .RN(n5), .Q(
        n66) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  SDFFRQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRQX2 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up2[1]) );
  SDFFRQX2 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n46), .CK(clk), .RN(n6), 
        .Q(up2[2]) );
  SDFFRQX4 up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n52), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  BUFX4 U3 ( .A(b1[1]), .Y(n4) );
  CLKBUFX1TH U4 ( .A(rst), .Y(n6) );
  CLKBUFX4TH U5 ( .A(rst), .Y(n5) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(up1[2]) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRX4 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n54), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRX4 up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(n55) );
  SDFFRX4 up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n53), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRHQX8 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n53), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  DLY1X1TH U38 ( .A(n47), .Y(n44) );
  DLY1X1TH U39 ( .A(n66), .Y(up1[0]) );
  INVXLTH U40 ( .A(n47), .Y(n46) );
  DLY1X1TH U41 ( .A(n51), .Y(n47) );
  INVXLTH U42 ( .A(n47), .Y(n48) );
  INVXLTH U43 ( .A(n51), .Y(n49) );
  DLY1X1TH U44 ( .A(test_se), .Y(n50) );
  INVXLTH U45 ( .A(test_se), .Y(n51) );
  INVXLTH U46 ( .A(n44), .Y(n52) );
  INVXLTH U47 ( .A(n44), .Y(n53) );
  INVXLTH U48 ( .A(n47), .Y(n54) );
  DLY1X1TH U49 ( .A(n55), .Y(up3[3]) );
  DLY1X1TH U50 ( .A(n67), .Y(up3[4]) );
endmodule


module sm_tc_91 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n21, n25, n26, n29;

  INVX4 U2 ( .A(n21), .Y(n25) );
  BUFX10 U3 ( .A(in[4]), .Y(n21) );
  OAI2BB2X2TH U4 ( .B0(n25), .B1(n6), .A0N(n29), .A1N(n25), .Y(out[1]) );
  NOR2X4 U5 ( .A(n29), .B(in[0]), .Y(n8) );
  CLKNAND2X2TH U6 ( .A(n8), .B(n26), .Y(n7) );
  INVX2TH U7 ( .A(in[2]), .Y(n26) );
  XNOR2X2TH U8 ( .A(n26), .B(n8), .Y(n5) );
  CLKBUFX1TH U9 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX2TH U10 ( .A(in[0]), .Y(out[0]) );
  NOR2BXLTH U11 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI22X2TH U12 ( .A0(n21), .A1(n26), .B0(n5), .B1(n25), .Y(out[2]) );
  OAI2BB2XLTH U13 ( .B0(n25), .B1(n4), .A0N(in[3]), .A1N(n25), .Y(out[3]) );
  XNOR2X4 U14 ( .A(n7), .B(in[3]), .Y(n4) );
  AO21X4 U15 ( .A0(in[0]), .A1(n29), .B0(n8), .Y(n6) );
  AOI31X2TH U16 ( .A0(n3), .A1(n4), .A2(n5), .B0(n25), .Y(out[4]) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX40 U18 ( .A(in[1]), .Y(n29) );
endmodule


module sm_tc_90 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n30, n31, n32, n36, n37;

  OR2X2 U2 ( .A(n36), .B(n5), .Y(n32) );
  BUFX10 U3 ( .A(in[1]), .Y(n30) );
  AO21X4 U4 ( .A0(in[0]), .A1(n30), .B0(n8), .Y(n6) );
  NOR2X6 U5 ( .A(n30), .B(in[0]), .Y(n8) );
  OAI2BB2XLTH U6 ( .B0(n36), .B1(n4), .A0N(in[3]), .A1N(n36), .Y(out[3]) );
  XNOR2X2TH U7 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2XL U8 ( .B0(n36), .B1(n6), .A0N(n30), .A1N(n36), .Y(out[1]) );
  INVX6 U9 ( .A(in[4]), .Y(n36) );
  NAND2XLTH U10 ( .A(n8), .B(n37), .Y(n7) );
  INVX2 U11 ( .A(in[2]), .Y(n37) );
  XNOR2X2TH U12 ( .A(n37), .B(n8), .Y(n5) );
  AOI31X2TH U13 ( .A0(n3), .A1(n4), .A2(n5), .B0(n36), .Y(out[4]) );
  OR2XLTH U14 ( .A(in[4]), .B(n37), .Y(n31) );
  NAND2X1TH U15 ( .A(n31), .B(n32), .Y(out[2]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U18 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U19 ( .A(out[4]), .Y(out[6]) );
endmodule


module sm_tc_89 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n18, n19, n23, n24;

  OAI22X1 U2 ( .A0(n18), .A1(n24), .B0(n23), .B1(n5), .Y(out[2]) );
  BUFX10 U3 ( .A(in[0]), .Y(n17) );
  OAI2BB2X4 U4 ( .B0(n23), .B1(n4), .A0N(in[3]), .A1N(n23), .Y(out[3]) );
  XNOR2X4 U5 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX16 U6 ( .A(n18), .Y(n23) );
  BUFX10 U7 ( .A(in[4]), .Y(n18) );
  INVX2TH U8 ( .A(in[2]), .Y(n24) );
  BUFX2 U9 ( .A(in[1]), .Y(n19) );
  OAI2BB2X1 U10 ( .B0(n23), .B1(n6), .A0N(n19), .A1N(n23), .Y(out[1]) );
  XNOR2X2TH U11 ( .A(n24), .B(n8), .Y(n5) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[6]) );
  AOI31X2TH U14 ( .A0(n3), .A1(n4), .A2(n5), .B0(n23), .Y(out[4]) );
  CLKBUFX1TH U15 ( .A(n17), .Y(out[0]) );
  AO21X2 U16 ( .A0(n17), .A1(n19), .B0(n8), .Y(n6) );
  NOR2X6 U17 ( .A(n19), .B(n17), .Y(n8) );
  NAND2XLTH U18 ( .A(n8), .B(n24), .Y(n7) );
  NOR2BXLTH U19 ( .AN(n6), .B(n17), .Y(n3) );
endmodule


module sm_tc_88 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  OAI2BB2X2 U5 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  XNOR2X1 U2 ( .A(n21), .B(n8), .Y(n5) );
  NOR2X4TH U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI22X1TH U4 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  XNOR2X1 U6 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKNAND2X2TH U7 ( .A(n8), .B(n21), .Y(n7) );
  CLKINVX2TH U8 ( .A(in[4]), .Y(n22) );
  CLKBUFX1TH U9 ( .A(in[0]), .Y(out[0]) );
  AO21XLTH U10 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n21) );
  OAI2BB2X1TH U12 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  INVXLTH U13 ( .A(out[4]), .Y(n18) );
  AOI31X2TH U14 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U16 ( .A(n18), .Y(out[5]) );
  INVXLTH U17 ( .A(n18), .Y(out[6]) );
endmodule


module add_22_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_22_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_22_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKAND2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_22_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_22_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X2 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_22_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n3, n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(n3) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKBUFX40 U3 ( .A(n3), .Y(SUM[1]) );
endmodule


module add_22 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  add_22_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n27, temp1_2_, 
        temp1_1_, temp1_0_}), .B({n29, in2[5:4], n16, n20, n19, in2[0]}), 
        .SUM(out3) );
  add_22_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, n17, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_22_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n27, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in3[6:4], n18, n26, n24, in3[0]}), .SUM(out2) );
  add_22_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n27, temp1_2_, 
        temp1_1_, temp1_0_}), .B({temp2_6_, n23, n17, n22, temp2_2_, temp2_1_, 
        temp2_0_}), .SUM(out) );
  add_22_DW01_add_4 add_30 ( .A({n28, in2[5:4], n16, n20, n19, in2[0]}), .B({
        in3[6:4], n18, n26, n24, in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_22_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX4 U1 ( .A(in2[3]), .Y(n16) );
  CLKINVX4 U2 ( .A(in3[2]), .Y(n25) );
  CLKBUFX2TH U3 ( .A(in3[3]), .Y(n18) );
  CLKBUFX2TH U4 ( .A(temp2_4_), .Y(n17) );
  BUFX2 U5 ( .A(in2[2]), .Y(n20) );
  BUFX2 U6 ( .A(in2[1]), .Y(n19) );
  CLKINVX1 U13 ( .A(temp2_3_), .Y(n21) );
  CLKBUFX2TH U14 ( .A(in3[1]), .Y(n24) );
  INVXLTH U15 ( .A(n21), .Y(n22) );
  CLKBUFX1TH U16 ( .A(temp2_5_), .Y(n23) );
  INVX1TH U17 ( .A(n25), .Y(n26) );
  CLKBUFX40 U18 ( .A(temp1_3_), .Y(n27) );
  DLY1X1TH U19 ( .A(in2[6]), .Y(n28) );
  DLY1X1TH U20 ( .A(in2[6]), .Y(n29) );
endmodule


module tc_sm_91 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(in[6]), .Y(n26) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n28) );
  INVXLTH U12 ( .A(in[5]), .Y(n27) );
  OAI21XLTH U13 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  CLKINVX1TH U14 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_90 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n21, n22, n23, n24, n25, n26, n28,
         n29, n30, n31, n32, n33;

  OR2X2 U3 ( .A(n28), .B(n10), .Y(n21) );
  OAI2BB1X4 U4 ( .A0N(n31), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI211XL U5 ( .A0(in[6]), .A1(n31), .B0(n7), .C0(n26), .Y(out[3]) );
  INVX2 U6 ( .A(n26), .Y(n25) );
  OR3XLTH U7 ( .A(n23), .B(n24), .C(n25), .Y(out[1]) );
  NAND3XL U8 ( .A(n21), .B(n22), .C(n26), .Y(out[2]) );
  OR2XLTH U9 ( .A(in[6]), .B(n32), .Y(n22) );
  INVXL U10 ( .A(in[6]), .Y(n28) );
  NOR2X2TH U11 ( .A(n28), .B(n12), .Y(n23) );
  NOR2XL U12 ( .A(in[6]), .B(n33), .Y(n24) );
  XNOR2X1TH U13 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVX2TH U14 ( .A(in[4]), .Y(n30) );
  CLKINVX1TH U15 ( .A(in[3]), .Y(n31) );
  NOR3X1TH U16 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U17 ( .A(in[1]), .Y(n33) );
  XNOR2XLTH U18 ( .A(n32), .B(n11), .Y(n10) );
  NOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI21XLTH U20 ( .A0(n9), .A1(n31), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U21 ( .A(in[6]), .Y(out[4]) );
  BUFX10 U22 ( .A(n8), .Y(n26) );
  NAND2BXLTH U23 ( .AN(in[0]), .B(n26), .Y(out[0]) );
  INVX2 U24 ( .A(in[5]), .Y(n29) );
  INVXLTH U25 ( .A(in[2]), .Y(n32) );
  OAI33X4 U26 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n29), .B2(
        n30), .Y(n8) );
endmodule


module tc_sm_89 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n9, n10, n11, n12, n18, n19, n20, n21, n22, n23, n25, n26, n27,
         n28;

  OAI211XL U3 ( .A0(in[6]), .A1(n21), .B0(n7), .C0(n28), .Y(out[3]) );
  OAI221XL U5 ( .A0(n18), .A1(n10), .B0(in[6]), .B1(n22), .C0(n28), .Y(out[2])
         );
  OAI221XL U6 ( .A0(n18), .A1(n12), .B0(in[6]), .B1(n23), .C0(n28), .Y(out[1])
         );
  CLKINVX1TH U7 ( .A(in[3]), .Y(n21) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U9 ( .A(in[6]), .Y(n18) );
  OAI21XLTH U10 ( .A0(n9), .A1(n21), .B0(in[6]), .Y(n7) );
  XNOR2XLTH U11 ( .A(n22), .B(n11), .Y(n10) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U13 ( .A(in[2]), .Y(n22) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U15 ( .A(in[1]), .Y(n23) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n28), .Y(out[0]) );
  INVX2 U18 ( .A(in[5]), .Y(n19) );
  INVXL U20 ( .A(in[4]), .Y(n20) );
  AOI33X4 U4 ( .A0(n20), .A1(n26), .A2(n19), .B0(n27), .B1(in[5]), .B2(in[4]), 
        .Y(n25) );
  CLKINVX40 U19 ( .A(in[6]), .Y(n26) );
  AOI21BX4 U21 ( .A0(n21), .A1(n9), .B0N(in[6]), .Y(n27) );
  CLKINVX40 U22 ( .A(n25), .Y(n28) );
endmodule


module tc_sm_88 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n28, n30, n31, n32, n33,
         n35, n36;

  CLKNAND2X8 U3 ( .A(n7), .B(n8), .Y(n11) );
  NAND3X4TH U4 ( .A(in[5]), .B(n35), .C(n14), .Y(n8) );
  NAND2X2 U5 ( .A(n6), .B(n5), .Y(out[3]) );
  OAI31XL U6 ( .A0(n8), .A1(n9), .A2(n31), .B0(in[6]), .Y(n5) );
  INVX4TH U7 ( .A(in[6]), .Y(n30) );
  AND2XLTH U9 ( .A(n9), .B(n31), .Y(n28) );
  NOR2X6 U10 ( .A(n28), .B(n30), .Y(n14) );
  INVXLTH U11 ( .A(in[3]), .Y(n31) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  OAI21XLTH U13 ( .A0(in[3]), .A1(n7), .B0(n30), .Y(n6) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n11), .Y(out[0]) );
  OAI221XLTH U16 ( .A0(n30), .A1(n13), .B0(in[6]), .B1(n33), .C0(n11), .Y(
        out[1]) );
  INVXLTH U17 ( .A(in[1]), .Y(n33) );
  XNOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n13) );
  OAI221XLTH U19 ( .A0(n30), .A1(n10), .B0(in[6]), .B1(n32), .C0(n11), .Y(
        out[2]) );
  XNOR2XLTH U20 ( .A(n32), .B(n12), .Y(n10) );
  NOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U22 ( .A(in[2]), .Y(n32) );
  INVXLTH U8 ( .A(n36), .Y(n35) );
  NAND3BX4 U23 ( .AN(in[5]), .B(n30), .C(n36), .Y(n7) );
  CLKINVX40 U24 ( .A(in[4]), .Y(n36) );
endmodule


module total_3_test_25 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n5, n6, n7, n8, n9, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_91 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_90 sm_tc_2 ( .out(b1), .in({n5, b[3:0]}) );
  sm_tc_89 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_88 sm_tc_4 ( .out(in1), .in(in) );
  add_22 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_91 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_90 tc_sm_2 ( .out(w6), .in({n7, w66[5:0]}) );
  tc_sm_89 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_88 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n54), .CK(clk), .RN(n9), .Q(
        up1[0]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n47), .CK(clk), .RN(n9), .Q(
        h) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n54), .CK(clk), .RN(n8), 
        .Q(up3[2]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n46), .CK(clk), .RN(n9), 
        .Q(up1[3]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n47), .CK(clk), .RN(n8), 
        .Q(up2[2]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n53), .CK(clk), .RN(n8), 
        .Q(up3[0]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n53), .CK(clk), .RN(n8), 
        .Q(up3[4]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n56), .CK(clk), .RN(n8), 
        .Q(up2[0]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n46), .CK(clk), .RN(n8), 
        .Q(up1[2]) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n55), .CK(clk), .RN(n8), 
        .Q(up2[4]) );
  SDFFRQXLTH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n50), .CK(clk), .RN(n8), 
        .Q(up2[1]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n56), .CK(clk), .RN(n8), 
        .Q(up3[1]) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n55), .CK(clk), .RN(n8), 
        .Q(up1[4]) );
  SDFFRQXLTH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n51), .CK(clk), .RN(n8), 
        .Q(up1[1]) );
  SDFFRQX2 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n50), .CK(clk), .RN(n8), 
        .Q(up2[3]) );
  BUFX2 U3 ( .A(b[4]), .Y(n5) );
  INVX12 U4 ( .A(n6), .Y(n7) );
  CLKBUFX4TH U5 ( .A(rst), .Y(n8) );
  CLKBUFX1TH U6 ( .A(rst), .Y(n9) );
  INVX2 U7 ( .A(w66[6]), .Y(n6) );
  SDFFRX4 up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n51), .CK(clk), .RN(n8), 
        .Q(up3[3]) );
  INVXLTH U40 ( .A(n49), .Y(n46) );
  INVXLTH U41 ( .A(n48), .Y(n47) );
  DLY1X1TH U42 ( .A(n52), .Y(n48) );
  DLY1X1TH U43 ( .A(n52), .Y(n49) );
  INVXLTH U44 ( .A(n49), .Y(n50) );
  INVXLTH U45 ( .A(n48), .Y(n51) );
  INVXLTH U46 ( .A(test_se), .Y(n52) );
  INVXLTH U47 ( .A(n49), .Y(n53) );
  INVXLTH U48 ( .A(n48), .Y(n54) );
  INVXLTH U49 ( .A(n49), .Y(n55) );
  INVXLTH U50 ( .A(n48), .Y(n56) );
endmodule


module sm_tc_87 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n21, n22, n23, n24, n25, n26, n30, n31, n34;

  NAND3XL U2 ( .A(n3), .B(n5), .C(n4), .Y(n25) );
  NOR2BXL U3 ( .AN(n6), .B(in[0]), .Y(n3) );
  XNOR2X2 U4 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKNAND2X2TH U6 ( .A(n21), .B(n22), .Y(n24) );
  AO21X1TH U7 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  INVX4 U8 ( .A(in[4]), .Y(n30) );
  BUFX2TH U9 ( .A(out[4]), .Y(out[5]) );
  INVX4 U10 ( .A(in[2]), .Y(n31) );
  AND2X1TH U11 ( .A(n25), .B(n26), .Y(out[4]) );
  OAI2BB2X4TH U12 ( .B0(n30), .B1(n6), .A0N(in[1]), .A1N(n30), .Y(out[1]) );
  BUFX2TH U13 ( .A(in[0]), .Y(out[0]) );
  NOR2X6 U14 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVXLTH U15 ( .A(n31), .Y(n21) );
  OAI2BB2XLTH U17 ( .B0(n4), .B1(n30), .A0N(in[3]), .A1N(n30), .Y(out[3]) );
  NAND2X2 U18 ( .A(n31), .B(n8), .Y(n23) );
  CLKINVX1TH U19 ( .A(n8), .Y(n22) );
  CLKBUFX1TH U20 ( .A(out[4]), .Y(out[6]) );
  INVXLTH U21 ( .A(n30), .Y(n26) );
  NAND2XLTH U22 ( .A(n8), .B(n31), .Y(n7) );
  OAI2BB2X2 U5 ( .B0(n30), .B1(n5), .A0N(n30), .A1N(in[2]), .Y(out[2]) );
  AND2X8 U16 ( .A(n23), .B(n24), .Y(n34) );
  CLKINVX40 U23 ( .A(n34), .Y(n5) );
endmodule


module sm_tc_86 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n4, n5, n6, n7, n8, n9, n20, n21, n22, n26, n27, n29, n30, n31, n32;

  AOI31X1 U2 ( .A0(n4), .A1(n5), .A2(n6), .B0(n32), .Y(out[4]) );
  OAI2BB2X2 U3 ( .B0(n32), .B1(n7), .A0N(in[1]), .A1N(n32), .Y(out[1]) );
  INVX2 U4 ( .A(in[4]), .Y(n27) );
  INVX1TH U5 ( .A(in[2]), .Y(n26) );
  NOR2X4 U6 ( .A(in[1]), .B(in[0]), .Y(n9) );
  XNOR2X4 U7 ( .A(n8), .B(in[3]), .Y(n5) );
  CLKBUFX1TH U8 ( .A(in[0]), .Y(out[0]) );
  OAI22X1TH U9 ( .A0(in[4]), .A1(n30), .B0(n32), .B1(n6), .Y(out[2]) );
  AO21XL U10 ( .A0(in[0]), .A1(in[1]), .B0(n9), .Y(n7) );
  CLKNAND2X2 U11 ( .A(n21), .B(n22), .Y(n6) );
  NAND2XLTH U12 ( .A(n9), .B(n30), .Y(n8) );
  NAND2XLTH U14 ( .A(n30), .B(n9), .Y(n21) );
  INVXLTH U15 ( .A(n9), .Y(n20) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X1TH U17 ( .B0(n32), .B1(n5), .A0N(in[3]), .A1N(n32), .Y(out[3]) );
  NOR2BXLTH U18 ( .AN(n7), .B(in[0]), .Y(n4) );
  CLKBUFX1TH U19 ( .A(out[4]), .Y(out[5]) );
  CLKINVX40 U13 ( .A(n26), .Y(n29) );
  CLKINVX40 U20 ( .A(n29), .Y(n30) );
  CLKINVX40 U21 ( .A(n27), .Y(n31) );
  CLKINVX40 U22 ( .A(n31), .Y(n32) );
  NAND2BX8 U23 ( .AN(n30), .B(n20), .Y(n22) );
endmodule


module sm_tc_85 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n27, n28, n29, n31, n34, n35, n38, n39, n40,
         n41;

  INVX2 U2 ( .A(out[4]), .Y(n31) );
  AOI31X2TH U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n35), .Y(out[4]) );
  CLKNAND2X4 U4 ( .A(n28), .B(n29), .Y(n4) );
  CLKNAND2X2 U6 ( .A(n7), .B(in[3]), .Y(n28) );
  CLKNAND2X4 U7 ( .A(n39), .B(n27), .Y(n29) );
  INVX1 U9 ( .A(in[3]), .Y(n27) );
  NOR2BXL U10 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVX6TH U11 ( .A(in[4]), .Y(n35) );
  OAI2BB2X1TH U13 ( .B0(n4), .B1(n35), .A0N(in[3]), .A1N(n35), .Y(out[3]) );
  OAI22X1TH U14 ( .A0(in[4]), .A1(n34), .B0(n35), .B1(n5), .Y(out[2]) );
  CLKBUFX1TH U15 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U16 ( .A(n31), .Y(out[6]) );
  NOR2X6 U17 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U18 ( .A(n31), .Y(out[5]) );
  INVX2 U20 ( .A(in[2]), .Y(n34) );
  XOR2X1 U5 ( .A(n34), .B(n38), .Y(n5) );
  CLKINVX40 U8 ( .A(n8), .Y(n38) );
  AO2B2X4 U12 ( .B0(in[4]), .B1(n40), .A0(in[1]), .A1N(in[4]), .Y(out[1]) );
  AND2X8 U19 ( .A(n8), .B(n34), .Y(n39) );
  CLKINVX40 U21 ( .A(n39), .Y(n7) );
  AOI21BX4 U22 ( .A0(in[0]), .A1(in[1]), .B0N(n41), .Y(n40) );
  CLKINVX40 U23 ( .A(n40), .Y(n6) );
  CLKINVX40 U24 ( .A(n8), .Y(n41) );
endmodule


module sm_tc_84 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n24, n25;

  BUFX2 U2 ( .A(out[4]), .Y(out[5]) );
  NOR2X2 U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X1 U4 ( .A(n7), .B(in[3]), .Y(n4) );
  AOI31X1 U5 ( .A0(n3), .A1(n4), .A2(n5), .B0(n24), .Y(out[4]) );
  XNOR2X1TH U6 ( .A(n25), .B(n8), .Y(n5) );
  CLKBUFX1TH U7 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X1 U8 ( .B0(n24), .B1(n4), .A0N(in[3]), .A1N(n24), .Y(out[3]) );
  CLKINVX2TH U9 ( .A(in[4]), .Y(n24) );
  CLKINVX1TH U10 ( .A(in[2]), .Y(n25) );
  OAI22X1TH U11 ( .A0(in[4]), .A1(n25), .B0(n24), .B1(n5), .Y(out[2]) );
  NAND2XLTH U12 ( .A(n8), .B(n25), .Y(n7) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2XL U15 ( .B0(n24), .B1(n6), .A0N(in[1]), .A1N(n24), .Y(out[1]) );
  AO21XLTH U16 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_21_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CLKXOR2X12 U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  CLKXOR2X2TH U2 ( .A(B[6]), .B(A[6]), .Y(n2) );
  AND2XLTH U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_21_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_21_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_21_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_21_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_21_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [6:2] carry;

  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  NAND2X2 U1 ( .A(B[5]), .B(n7), .Y(n8) );
  NAND2X3 U2 ( .A(n6), .B(A[5]), .Y(n9) );
  CLKNAND2X4 U3 ( .A(n8), .B(n9), .Y(n2) );
  CLKINVX3 U4 ( .A(B[5]), .Y(n6) );
  INVXL U5 ( .A(A[5]), .Y(n7) );
  XOR2X3 U6 ( .A(n2), .B(n10), .Y(SUM[5]) );
  CLKXOR2X2TH U7 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U8 ( .A(B[0]), .B(A[0]), .Y(n1) );
  NAND2XLTH U9 ( .A(A[5]), .B(B[5]), .Y(n5) );
  NAND2XLTH U10 ( .A(n10), .B(B[5]), .Y(n4) );
  NAND2XLTH U11 ( .A(n10), .B(A[5]), .Y(n3) );
  NAND3X2 U12 ( .A(n3), .B(n4), .C(n5), .Y(carry[6]) );
  CLKBUFX40 U13 ( .A(carry[5]), .Y(n10) );
endmodule


module add_21 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n18, n19, n20, n21, n22, n23, n24, n25, n26;

  add_21_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n25, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in2[6:5], n23, in2[3], n19, n26, in2[0]}), 
        .SUM(out3) );
  add_21_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B({in[6:5], n22, in[3:0]}), .SUM(out1) );
  add_21_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n25, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in3[6:3], n24, n18, in3[0]}), .SUM(out2) );
  add_21_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n25, temp1_2_, 
        temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_21_DW01_add_4 add_30 ( .A({in2[6:5], n23, in2[3], n19, n26, in2[0]}), 
        .B({in3[6:3], n24, in3[1:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_21_DW01_add_5 add_29 ( .A({in[6:5], n21, in[3:0]}), .B(in1), .SUM({
        temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_})
         );
  BUFX2 U1 ( .A(in3[1]), .Y(n18) );
  INVX2 U2 ( .A(in[4]), .Y(n20) );
  BUFX2 U3 ( .A(in2[2]), .Y(n19) );
  CLKBUFX1TH U4 ( .A(in2[4]), .Y(n23) );
  INVXLTH U5 ( .A(n20), .Y(n21) );
  INVXLTH U6 ( .A(n20), .Y(n22) );
  CLKBUFX40 U13 ( .A(in3[2]), .Y(n24) );
  CLKBUFX40 U14 ( .A(temp1_3_), .Y(n25) );
  CLKBUFX40 U15 ( .A(in2[1]), .Y(n26) );
endmodule


module tc_sm_87 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U10 ( .A(in[4]), .Y(n28) );
  INVXLTH U11 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_86 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n11, n12, n25, n26, n27, n29, n30, n31, n32, n33, n34,
         n36, n37, n38, n39, n40;

  INVXLTH U3 ( .A(in[4]), .Y(n31) );
  INVX4 U4 ( .A(n27), .Y(out[4]) );
  INVX2 U5 ( .A(in[6]), .Y(n27) );
  AOI33X4 U6 ( .A0(n31), .A1(n27), .A2(n30), .B0(n26), .B1(in[5]), .B2(in[4]), 
        .Y(n25) );
  CLKINVX32 U7 ( .A(n25), .Y(n8) );
  AOI21BX2TH U8 ( .A0(n32), .A1(n9), .B0N(in[6]), .Y(n26) );
  INVXL U10 ( .A(out[4]), .Y(n29) );
  OAI221X1 U11 ( .A0(n29), .A1(n12), .B0(out[4]), .B1(n34), .C0(n8), .Y(out[1]) );
  OAI211X2TH U12 ( .A0(out[4]), .A1(n32), .B0(n7), .C0(n8), .Y(out[3]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  CLKINVX1TH U15 ( .A(in[3]), .Y(n32) );
  NOR3X1TH U16 ( .A(in[1]), .B(n36), .C(in[0]), .Y(n9) );
  INVX2 U18 ( .A(in[5]), .Y(n30) );
  INVXLTH U19 ( .A(in[1]), .Y(n34) );
  XNOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U22 ( .A(n36), .Y(n33) );
  DLY1X1TH U9 ( .A(in[2]), .Y(n36) );
  AOI221X4 U13 ( .A0(out[4]), .A1(n39), .B0(n27), .B1(n36), .C0(n38), .Y(n37)
         );
  CLKINVX40 U17 ( .A(n37), .Y(out[2]) );
  CLKINVX40 U23 ( .A(n8), .Y(n38) );
  CLKXOR2X12 U24 ( .A(n33), .B(n11), .Y(n39) );
  OA21X4 U25 ( .A0(n9), .A1(n32), .B0(out[4]), .Y(n40) );
  CLKINVX40 U26 ( .A(n40), .Y(n7) );
endmodule


module tc_sm_85 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n11, n12, n13, n27, n28, n30, n31, n32, n33, n35,
         n36, n37, n38, n39, n40;

  CLKNAND2X2TH U4 ( .A(n5), .B(n6), .Y(out[3]) );
  OR2XLTH U5 ( .A(n30), .B(n13), .Y(n27) );
  OR2XLTH U6 ( .A(in[6]), .B(n33), .Y(n28) );
  NAND3XLTH U7 ( .A(n27), .B(n28), .C(n11), .Y(out[1]) );
  INVX2TH U8 ( .A(in[6]), .Y(n30) );
  OR3X1TH U9 ( .A(in[5]), .B(in[6]), .C(in[4]), .Y(n7) );
  OAI2B11X2TH U10 ( .A1N(n9), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n8) );
  OAI21XL U11 ( .A0(in[3]), .A1(n7), .B0(n30), .Y(n6) );
  OAI31XL U12 ( .A0(n8), .A1(n9), .A2(n31), .B0(in[6]), .Y(n5) );
  NOR3X1TH U13 ( .A(in[1]), .B(n36), .C(in[0]), .Y(n9) );
  INVXLTH U14 ( .A(in[1]), .Y(n33) );
  XNOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n13) );
  INVXLTH U17 ( .A(n36), .Y(n32) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U19 ( .A(in[3]), .Y(n31) );
  CLKBUFX1TH U20 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U22 ( .AN(in[0]), .B(n11), .Y(out[0]) );
  CLKBUFX40 U3 ( .A(n38), .Y(n35) );
  DLY1X1TH U16 ( .A(in[2]), .Y(n36) );
  OA21X4 U21 ( .A0(n30), .A1(n8), .B0(n7), .Y(n37) );
  CLKINVX40 U23 ( .A(n37), .Y(n11) );
  AOI221X4 U24 ( .A0(in[6]), .A1(n40), .B0(n30), .B1(n36), .C0(n39), .Y(n38)
         );
  CLKINVX40 U25 ( .A(n35), .Y(out[2]) );
  CLKINVX40 U26 ( .A(n11), .Y(n39) );
  CLKXOR2X12 U27 ( .A(n32), .B(n12), .Y(n40) );
endmodule


module tc_sm_84 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n22, n23, n24, n25, n27, n28,
         n29;

  OAI221XL U4 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[2])
         );
  OAI221XL U5 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[1])
         );
  OAI211XL U6 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
  INVXLTH U9 ( .A(in[6]), .Y(n20) );
  CLKINVX1TH U10 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U12 ( .A(in[4]), .Y(n22) );
  INVXLTH U13 ( .A(in[5]), .Y(n21) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U15 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U17 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U19 ( .A(in[2]), .Y(n24) );
  OAI21XLTH U20 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  NAND2BXLTH U21 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  AOI33X4 U3 ( .A0(n22), .A1(n28), .A2(n21), .B0(n29), .B1(in[5]), .B2(in[4]), 
        .Y(n27) );
  CLKINVX40 U7 ( .A(n27), .Y(n8) );
  CLKINVX40 U8 ( .A(in[6]), .Y(n28) );
  AOI21BX4 U22 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n29) );
endmodule


module total_3_test_26 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n5, n6, n7, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_87 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_86 sm_tc_2 ( .out(b1), .in({b[4:1], n5}) );
  sm_tc_85 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_84 sm_tc_4 ( .out(in1), .in(in) );
  add_21 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_87 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_86 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_85 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_84 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up3[3]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n59), .CK(clk), .RN(n6), 
        .Q(up3[2]) );
  SDFFRQXL up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n57), .CK(clk), .RN(n6), 
        .Q(up1[1]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n55), .CK(clk), .RN(n7), .Q(
        h) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up2[4]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n58), .CK(clk), .RN(n6), 
        .Q(up2[3]) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n57), .CK(clk), .RN(n7), 
        .Q(up1[4]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n55), .CK(clk), .RN(n6), 
        .Q(up3[0]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up1[3]) );
  SDFFRQX1TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n59), .CK(clk), .RN(n6), 
        .Q(up3[4]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n55), .CK(clk), .RN(n6), 
        .Q(up2[0]) );
  SDFFRHQX2 up1_reg_2_ ( .D(w6[2]), .SI(n61), .SE(n55), .CK(clk), .RN(n6), .Q(
        up1[2]) );
  CLKBUFX4 U3 ( .A(b[0]), .Y(n5) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n6) );
  CLKBUFX1TH U5 ( .A(rst), .Y(n7) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up2[1]) );
  SDFFRX4 up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n58), .CK(clk), .RN(n6), .Q(
        up1[0]) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up3[1]) );
  SDFFRX4 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n50), .CK(clk), .RN(n7), 
        .Q(up2[2]) );
  DLY1X1TH U38 ( .A(n53), .Y(n50) );
  DLY1X1TH U39 ( .A(n54), .Y(n51) );
  DLY1X1TH U40 ( .A(n56), .Y(n52) );
  INVXLTH U41 ( .A(n52), .Y(n53) );
  INVXLTH U42 ( .A(n56), .Y(n54) );
  DLY1X1TH U43 ( .A(test_se), .Y(n55) );
  INVXLTH U44 ( .A(test_se), .Y(n56) );
  INVXLTH U45 ( .A(n52), .Y(n57) );
  INVXLTH U46 ( .A(n52), .Y(n58) );
  INVXLTH U47 ( .A(n52), .Y(n59) );
  INVXLTH U48 ( .A(up1[1]), .Y(n60) );
  INVXLTH U49 ( .A(n60), .Y(n61) );
endmodule


module sm_tc_83 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n21, n25, n26, n29, n30;

  OAI22X1 U3 ( .A0(n21), .A1(n29), .B0(n25), .B1(n5), .Y(out[2]) );
  XNOR2X2 U4 ( .A(n29), .B(n8), .Y(n5) );
  BUFX2 U5 ( .A(in[4]), .Y(n21) );
  INVX1TH U6 ( .A(in[2]), .Y(n26) );
  CLKBUFX1TH U7 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X2 U8 ( .B0(n25), .B1(n6), .A0N(in[1]), .A1N(n25), .Y(out[1]) );
  AO21X2 U9 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X6 U10 ( .A(in[1]), .B(in[0]), .Y(n8) );
  BUFX2 U11 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2X1 U12 ( .B0(n25), .B1(n4), .A0N(in[3]), .A1N(n25), .Y(out[3]) );
  CLKBUFX1TH U13 ( .A(in[0]), .Y(out[0]) );
  AOI31X2TH U15 ( .A0(n3), .A1(n4), .A2(n5), .B0(n25), .Y(out[4]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVX4 U17 ( .A(n21), .Y(n25) );
  CLKBUFX40 U2 ( .A(n26), .Y(n29) );
  XOR2X1 U14 ( .A(n30), .B(in[3]), .Y(n4) );
  CLKAND2X12 U18 ( .A(n8), .B(n29), .Y(n30) );
endmodule


module sm_tc_82 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n19, n20, n21, n22, n23, n24, n25, n29, n30,
         n33, n34;

  NAND2XL U2 ( .A(n8), .B(n30), .Y(n7) );
  NOR2X6 U3 ( .A(n34), .B(in[0]), .Y(n8) );
  CLKNAND2X2 U4 ( .A(n20), .B(n21), .Y(n5) );
  OAI2BB2X2 U5 ( .B0(n29), .B1(n6), .A0N(n34), .A1N(n29), .Y(out[1]) );
  INVX2 U6 ( .A(in[4]), .Y(n29) );
  OAI22X2 U7 ( .A0(in[4]), .A1(n30), .B0(n29), .B1(n5), .Y(out[2]) );
  NAND2XLTH U8 ( .A(n30), .B(n8), .Y(n20) );
  INVX2 U9 ( .A(in[2]), .Y(n30) );
  AO21XLTH U10 ( .A0(in[0]), .A1(n34), .B0(n8), .Y(n6) );
  AOI31X4TH U11 ( .A0(n3), .A1(n4), .A2(n5), .B0(n29), .Y(out[4]) );
  NAND2X4TH U12 ( .A(n24), .B(n25), .Y(n4) );
  CLKNAND2X4TH U13 ( .A(n22), .B(n23), .Y(n25) );
  OAI2BB2X2TH U15 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  INVXLTH U16 ( .A(in[3]), .Y(n23) );
  INVXLTH U17 ( .A(n7), .Y(n22) );
  NAND2XLTH U18 ( .A(n7), .B(in[3]), .Y(n24) );
  INVXLTH U19 ( .A(n8), .Y(n19) );
  NOR2BXLTH U20 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U21 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U22 ( .A(out[4]), .Y(out[6]) );
  BUFX2TH U23 ( .A(in[0]), .Y(out[0]) );
  AND2X8 U14 ( .A(in[2]), .B(n19), .Y(n33) );
  CLKINVX40 U24 ( .A(n33), .Y(n21) );
  CLKBUFX40 U25 ( .A(in[1]), .Y(n34) );
endmodule


module sm_tc_81 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n20, n21, n23, n33, n26, n27, n30, n32;

  OAI2BB2X1 U2 ( .B0(n27), .B1(n6), .A0N(n32), .A1N(n27), .Y(out[1]) );
  OAI22X2 U3 ( .A0(n20), .A1(n26), .B0(n27), .B1(n5), .Y(out[2]) );
  OAI2BB2X4 U4 ( .B0(n27), .B1(n4), .A0N(in[3]), .A1N(n27), .Y(out[3]) );
  INVX4 U5 ( .A(n20), .Y(n27) );
  INVX2TH U6 ( .A(in[2]), .Y(n26) );
  BUFX8 U8 ( .A(in[4]), .Y(n20) );
  XNOR2X1 U9 ( .A(n26), .B(n8), .Y(n5) );
  NOR2X4 U10 ( .A(n32), .B(in[0]), .Y(n8) );
  XNOR2X1TH U11 ( .A(n7), .B(in[3]), .Y(n4) );
  AND2X6 U12 ( .A(n21), .B(n20), .Y(out[4]) );
  INVXLTH U13 ( .A(out[4]), .Y(n23) );
  NAND3X1 U14 ( .A(n3), .B(n4), .C(n5), .Y(n21) );
  CLKBUFX1TH U16 ( .A(in[0]), .Y(out[0]) );
  CLKINVX1TH U17 ( .A(n23), .Y(n33) );
  AO21X1 U18 ( .A0(in[0]), .A1(n32), .B0(n8), .Y(n6) );
  NOR2BXLTH U19 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U20 ( .A(n23), .Y(out[6]) );
  AND2X8 U7 ( .A(n8), .B(n26), .Y(n30) );
  CLKINVX40 U15 ( .A(n30), .Y(n7) );
  CLKBUFX40 U21 ( .A(n33), .Y(out[5]) );
  CLKBUFX40 U22 ( .A(in[1]), .Y(n32) );
endmodule


module sm_tc_80 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n18, n19, n20, n22, n25, n26;

  AOI31X2 U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n26), .Y(out[4]) );
  CLKNAND2X2 U3 ( .A(n17), .B(n18), .Y(n20) );
  NAND2X2 U4 ( .A(n7), .B(in[3]), .Y(n19) );
  NAND2X4 U5 ( .A(n19), .B(n20), .Y(n4) );
  CLKINVX2 U6 ( .A(n7), .Y(n17) );
  INVX2 U7 ( .A(in[3]), .Y(n18) );
  NAND2XL U8 ( .A(n8), .B(n25), .Y(n7) );
  OAI2BB2X1 U9 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  NOR2X3TH U10 ( .A(in[1]), .B(in[0]), .Y(n8) );
  NOR2BXLTH U11 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVX1TH U12 ( .A(out[4]), .Y(n22) );
  OAI2BB2X2TH U13 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n26), .Y(out[1]) );
  CLKBUFX1TH U14 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1 U15 ( .A(n25), .B(n8), .Y(n5) );
  CLKINVX2TH U16 ( .A(in[4]), .Y(n26) );
  CLKINVX1TH U17 ( .A(in[2]), .Y(n25) );
  INVXLTH U18 ( .A(n22), .Y(out[5]) );
  OAI22X1TH U19 ( .A0(in[4]), .A1(n25), .B0(n26), .B1(n5), .Y(out[2]) );
  INVXLTH U20 ( .A(n22), .Y(out[6]) );
  AO21XLTH U21 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_20_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3;
  wire   [6:2] carry;

  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(A[0]), .B(B[0]), .Y(n1) );
  CLKXOR2X8 U4 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  XNOR2X1 U3 ( .A(n3), .B(A[6]), .Y(n2) );
  CLKINVX40 U5 ( .A(B[6]), .Y(n3) );
endmodule


module add_20_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR2X4 U3 ( .A(A[6]), .B(B[6]), .Y(n2) );
  CLKXOR2X8 U4 ( .A(n3), .B(carry[6]), .Y(SUM[6]) );
  CLKINVX20 U5 ( .A(n2), .Y(n3) );
endmodule


module add_20_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_20_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_20_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [6:2] carry;

  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  INVX2 U1 ( .A(carry[4]), .Y(n7) );
  NAND3X2 U2 ( .A(n3), .B(n4), .C(n5), .Y(carry[5]) );
  CLKNAND2X4 U3 ( .A(n8), .B(n9), .Y(SUM[4]) );
  INVXLTH U5 ( .A(n2), .Y(n6) );
  CLKXOR2X4 U6 ( .A(A[4]), .B(B[4]), .Y(n2) );
  CLKXOR2X2TH U7 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  NAND2XLTH U8 ( .A(n6), .B(carry[4]), .Y(n9) );
  NAND2XLTH U9 ( .A(B[4]), .B(A[4]), .Y(n5) );
  NAND2XLTH U10 ( .A(carry[4]), .B(B[4]), .Y(n3) );
  NAND2XLTH U11 ( .A(carry[4]), .B(A[4]), .Y(n4) );
  AND2XLTH U12 ( .A(B[0]), .B(A[0]), .Y(n1) );
  AND2X8 U4 ( .A(n2), .B(n7), .Y(n10) );
  CLKINVX40 U13 ( .A(n10), .Y(n8) );
endmodule


module add_20_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR2X3TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_20 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23;

  add_20_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n20, temp1_2_, 
        n18, temp1_0_}), .B({n23, in2[5:3], n16, n21, in2[0]}), .SUM(out3) );
  add_20_DW01_add_1 add_33 ( .A({n19, temp2_5_, n15, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_20_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n20, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in3[6:2], n17, n14}), .SUM(out2) );
  add_20_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n20, temp1_2_, 
        n18, temp1_0_}), .B({n19, temp2_5_, n15, temp2_3_, temp2_2_, temp2_1_, 
        temp2_0_}), .SUM(out) );
  add_20_DW01_add_4 add_30 ( .A({n22, in2[5:3], n16, n21, in2[0]}), .B({
        in3[6:2], n17, in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}) );
  add_20_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX4 U1 ( .A(temp2_4_), .Y(n15) );
  CLKBUFX2 U2 ( .A(in2[2]), .Y(n16) );
  BUFX2 U3 ( .A(in3[0]), .Y(n14) );
  CLKBUFX2TH U4 ( .A(in3[1]), .Y(n17) );
  CLKBUFX40 U5 ( .A(temp1_1_), .Y(n18) );
  CLKBUFX40 U6 ( .A(temp2_6_), .Y(n19) );
  CLKBUFX40 U13 ( .A(temp1_3_), .Y(n20) );
  CLKBUFX40 U14 ( .A(in2[1]), .Y(n21) );
  DLY1X1TH U15 ( .A(in2[6]), .Y(n22) );
  DLY1X1TH U16 ( .A(in2[6]), .Y(n23) );
endmodule


module tc_sm_83 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U10 ( .A(in[4]), .Y(n28) );
  INVXLTH U11 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_82 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n17, n18, n20, n21, n22, n23, n24,
         n25, n27;

  OAI221X2TH U3 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n18), .Y(
        out[1]) );
  BUFX8 U4 ( .A(n8), .Y(n18) );
  OA21XL U5 ( .A0(in[6]), .A1(n23), .B0(n7), .Y(n17) );
  NAND2XLTH U6 ( .A(n17), .B(n18), .Y(out[3]) );
  INVXLTH U7 ( .A(in[6]), .Y(n20) );
  OAI221X1 U8 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n18), .Y(out[2])
         );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  OAI33X4 U10 ( .A0(in[4]), .A1(in[6]), .A2(n27), .B0(n13), .B1(n21), .B2(n22), 
        .Y(n8) );
  OAI2BB1X4 U11 ( .A0N(n23), .A1N(n9), .B0(in[6]), .Y(n13) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n23) );
  INVXLTH U13 ( .A(in[4]), .Y(n22) );
  INVXLTH U14 ( .A(n27), .Y(n21) );
  XNOR2XLTH U15 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U17 ( .A(in[2]), .Y(n24) );
  OAI21XLTH U18 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  INVXLTH U19 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U21 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  CLKBUFX1TH U22 ( .A(in[6]), .Y(out[4]) );
  CLKBUFX40 U23 ( .A(in[5]), .Y(n27) );
endmodule


module tc_sm_81 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n18, n19, n20, n21, n22, n24, n25, n26,
         n27, n28;

  INVX2 U3 ( .A(in[6]), .Y(n21) );
  INVX2 U4 ( .A(n20), .Y(n8) );
  OR2XLTH U5 ( .A(n21), .B(n12), .Y(n18) );
  OR2XLTH U6 ( .A(in[6]), .B(n28), .Y(n19) );
  NAND3XLTH U7 ( .A(n18), .B(n19), .C(n8), .Y(out[1]) );
  AOI33X2 U8 ( .A0(n25), .A1(n21), .A2(n24), .B0(n22), .B1(in[5]), .B2(in[4]), 
        .Y(n20) );
  AOI21BX2TH U9 ( .A0(n26), .A1(n9), .B0N(in[6]), .Y(n22) );
  INVXLTH U10 ( .A(in[4]), .Y(n25) );
  INVX2TH U11 ( .A(in[5]), .Y(n24) );
  OAI221XLTH U12 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n27), .C0(n8), .Y(
        out[2]) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n26) );
  NOR3X1TH U14 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U15 ( .A(in[1]), .Y(n28) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U17 ( .A(n27), .B(n11), .Y(n10) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U19 ( .A(in[2]), .Y(n27) );
  OAI21XLTH U20 ( .A0(n9), .A1(n26), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U21 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U22 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211XLTH U23 ( .A0(in[6]), .A1(n26), .B0(n7), .C0(n8), .Y(out[3]) );
endmodule


module tc_sm_80 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n9, n10, n11, n12, n19, n20, n22, n23, n24, n26, n27, n28, n29,
         n30, n31;

  OAI211XLTH U3 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n31), .Y(out[3]) );
  OAI221X1 U4 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n31), .Y(out[1])
         );
  INVX1TH U6 ( .A(in[5]), .Y(n20) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n22) );
  OAI221X1TH U9 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n31), .Y(
        out[2]) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U11 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U13 ( .A(in[2]), .Y(n23) );
  OAI21XLTH U14 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  INVXLTH U15 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U18 ( .A(in[6]), .Y(n19) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n31), .Y(out[0]) );
  DLY1X1TH U5 ( .A(in[4]), .Y(n26) );
  AOI33X4 U7 ( .A0(n28), .A1(n29), .A2(n20), .B0(n30), .B1(in[5]), .B2(in[4]), 
        .Y(n27) );
  CLKINVX40 U20 ( .A(n26), .Y(n28) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n29) );
  AOI21BX4 U22 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n30) );
  CLKINVX40 U23 ( .A(n27), .Y(n31) );
endmodule


module total_3_test_27 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n5, n6, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_83 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_82 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_81 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_80 sm_tc_4 ( .out(in1), .in(in) );
  add_20 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_83 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_82 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_81 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_80 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n52), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n50), .CK(clk), .RN(n5), .Q(
        up1[0]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n46), .CK(clk), .RN(n6), .Q(
        h) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n54), .CK(clk), .RN(n5), 
        .Q(up3[3]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n53), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRQX1TH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRQX2 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n52), .CK(clk), .RN(rst), 
        .Q(up2[1]) );
  SDFFRQX2 up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n54), .CK(clk), .RN(n5), 
        .Q(up3[4]) );
  SDFFRQX1TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQX2 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up1[3]) );
  BUFX3TH U3 ( .A(rst), .Y(n5) );
  CLKBUFX1TH U5 ( .A(rst), .Y(n6) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n53), .CK(clk), .RN(n5), 
        .Q(up1[2]) );
  SDFFRX4 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  SDFFRHQX8 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up2[2]) );
  DLY1X1TH U37 ( .A(n47), .Y(n45) );
  INVXLTH U38 ( .A(n47), .Y(n46) );
  DLY1X1TH U39 ( .A(n51), .Y(n47) );
  INVXLTH U40 ( .A(n47), .Y(n48) );
  INVXLTH U41 ( .A(n51), .Y(n49) );
  DLY1X1TH U42 ( .A(test_se), .Y(n50) );
  INVXLTH U43 ( .A(test_se), .Y(n51) );
  INVXLTH U44 ( .A(n45), .Y(n52) );
  INVXLTH U45 ( .A(n45), .Y(n53) );
  INVXLTH U46 ( .A(n47), .Y(n54) );
endmodule


module sm_tc_79 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n29, n3, n4, n5, n6, n7, n8, n21, n22, n25, n26, n27;

  NOR2X4 U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  NAND2X2 U3 ( .A(n8), .B(n21), .Y(n7) );
  CLKINVX1TH U5 ( .A(in[2]), .Y(n21) );
  CLKBUFX1TH U6 ( .A(out[4]), .Y(out[6]) );
  OAI22X4 U7 ( .A0(in[4]), .A1(n21), .B0(n27), .B1(n5), .Y(out[2]) );
  AOI31X1 U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n27), .Y(n29) );
  CLKBUFX1TH U9 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X4TH U10 ( .B0(n27), .B1(n6), .A0N(in[1]), .A1N(n27), .Y(out[1]) );
  XNOR2X1TH U11 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX2TH U12 ( .A(in[4]), .Y(n22) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  AO21XLTH U16 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  XNOR2X1 U4 ( .A(in[2]), .B(n25), .Y(n5) );
  CLKINVX40 U13 ( .A(n8), .Y(n25) );
  OAI2B2X2 U17 ( .A1N(in[3]), .A0(n26), .B0(n27), .B1(n4), .Y(out[3]) );
  CLKINVX40 U18 ( .A(n22), .Y(n26) );
  CLKINVX40 U19 ( .A(n26), .Y(n27) );
  CLKBUFX40 U20 ( .A(n29), .Y(out[4]) );
endmodule


module sm_tc_78 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n24, n28, n29, n31, n32;

  BUFX6 U2 ( .A(in[4]), .Y(n24) );
  OAI22X2TH U3 ( .A0(n24), .A1(n28), .B0(n29), .B1(n5), .Y(out[2]) );
  NOR2BXL U4 ( .AN(n6), .B(out[0]), .Y(n3) );
  BUFX4TH U6 ( .A(in[0]), .Y(out[0]) );
  INVX2 U7 ( .A(in[2]), .Y(n28) );
  AO21XLTH U10 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  XNOR2X4TH U11 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX2TH U12 ( .A(n24), .Y(n29) );
  AOI31X2TH U13 ( .A0(n3), .A1(n4), .A2(n5), .B0(n29), .Y(out[6]) );
  OAI2BB2XLTH U14 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  CLKBUFX1TH U15 ( .A(out[6]), .Y(out[5]) );
  CLKBUFX1TH U16 ( .A(out[6]), .Y(out[4]) );
  AO2B2BX4 U5 ( .A0(n24), .A1N(n6), .B0(in[1]), .B1N(n24), .Y(out[1]) );
  OR2X8 U8 ( .A(in[1]), .B(out[0]), .Y(n31) );
  CLKINVX40 U9 ( .A(n31), .Y(n8) );
  XOR2X1 U17 ( .A(n28), .B(n31), .Y(n5) );
  AND2X8 U18 ( .A(n8), .B(n28), .Y(n32) );
  CLKINVX40 U19 ( .A(n32), .Y(n7) );
endmodule


module sm_tc_77 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n32, n33, n35, n36, n37;

  INVX2 U2 ( .A(in[2]), .Y(n32) );
  XNOR2X1 U3 ( .A(n32), .B(n8), .Y(n5) );
  INVX2TH U4 ( .A(in[4]), .Y(n33) );
  NOR2BXLTH U5 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI22X2TH U6 ( .A0(in[4]), .A1(n32), .B0(n37), .B1(n5), .Y(out[2]) );
  AOI31X4 U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n37), .Y(out[6]) );
  XNOR2X2TH U8 ( .A(n7), .B(in[3]), .Y(n4) );
  AO21XLTH U10 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2X4 U11 ( .B0(n37), .B1(n6), .A0N(in[1]), .A1N(n37), .Y(out[1]) );
  CLKBUFX1TH U13 ( .A(out[6]), .Y(out[5]) );
  CLKBUFX1TH U14 ( .A(out[6]), .Y(out[4]) );
  BUFX2TH U15 ( .A(in[0]), .Y(out[0]) );
  NAND2XLTH U16 ( .A(n8), .B(n32), .Y(n7) );
  OAI2B2X2 U9 ( .A1N(in[3]), .A0(n36), .B0(n37), .B1(n4), .Y(out[3]) );
  OR2X8 U12 ( .A(in[1]), .B(in[0]), .Y(n35) );
  CLKINVX40 U17 ( .A(n35), .Y(n8) );
  CLKINVX40 U18 ( .A(n33), .Y(n36) );
  CLKINVX40 U19 ( .A(n36), .Y(n37) );
endmodule


module sm_tc_76 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  NOR2X2 U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X1TH U3 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U4 ( .A(n8), .B(n21), .Y(n7) );
  OAI2BB2X1TH U5 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  XNOR2X1TH U6 ( .A(n21), .B(n8), .Y(n5) );
  OAI2BB2X2TH U7 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  CLKBUFX1TH U8 ( .A(in[0]), .Y(out[0]) );
  OAI22X4TH U9 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  INVXLTH U10 ( .A(n18), .Y(out[6]) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n21) );
  CLKINVX2TH U12 ( .A(in[4]), .Y(n22) );
  INVXLTH U13 ( .A(out[4]), .Y(n18) );
  AOI31X2TH U14 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U16 ( .A(n18), .Y(out[5]) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_19_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_19_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_19_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_19_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR3X2 U3 ( .A(n3), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
  CLKINVX40 U5 ( .A(A[6]), .Y(n3) );
endmodule


module add_19_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHX2TH U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_19_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n3, n4, n5, n6, n7, n8;
  wire   [6:2] carry;

  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX4TH U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX2TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XNOR2X2TH U1 ( .A(n6), .B(n7), .Y(SUM[2]) );
  NAND2XLTH U2 ( .A(n7), .B(B[2]), .Y(n4) );
  XNOR2X4TH U3 ( .A(B[2]), .B(A[2]), .Y(n6) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X2TH U5 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2XLTH U7 ( .A(A[2]), .B(B[2]), .Y(n5) );
  NAND2XLTH U8 ( .A(n7), .B(A[2]), .Y(n3) );
  CLKBUFX40 U6 ( .A(carry[2]), .Y(n7) );
  AND3X8 U9 ( .A(n3), .B(n4), .C(n5), .Y(n8) );
  CLKINVX40 U10 ( .A(n8), .Y(carry[3]) );
endmodule


module add_19 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   n24, temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_,
         temp2_0_, temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_,
         temp1_0_, n18, n19, n20, n21, n23;

  add_19_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n20, 
        temp1_1_, temp1_0_}), .B({n21, in2[5:4], n19, in2[2:0]}), .SUM(out3)
         );
  add_19_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, n23, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .B(in), .SUM({n24, out1[5:0]}) );
  add_19_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n20, 
        temp1_1_, temp1_0_}), .B(in3), .SUM(out2) );
  add_19_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, n20, 
        temp1_1_, n18}), .B({temp2_6_, temp2_5_, n23, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_19_DW01_add_4 add_30 ( .A({n21, in2[5:4], n19, in2[2:0]}), .B(in3), 
        .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, 
        temp2_0_}) );
  add_19_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2 U1 ( .A(temp1_2_), .Y(n20) );
  CLKBUFX1TH U2 ( .A(in2[6]), .Y(n21) );
  CLKBUFX1TH U3 ( .A(temp1_0_), .Y(n18) );
  CLKBUFX1TH U4 ( .A(in2[3]), .Y(n19) );
  CLKBUFX40 U5 ( .A(n24), .Y(out1[6]) );
  CLKBUFX40 U6 ( .A(temp2_4_), .Y(n23) );
endmodule


module tc_sm_79 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U10 ( .A(in[4]), .Y(n28) );
  INVXLTH U11 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_78 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n23, n24, n25, n26, n28, n29;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OAI211XLTH U3 ( .A0(in[6]), .A1(n24), .B0(n5), .C0(n6), .Y(out[3]) );
  INVXLTH U4 ( .A(in[6]), .Y(n23) );
  NOR3X1TH U6 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U8 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U9 ( .A(in[2]), .Y(n25) );
  XOR2XLTH U10 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI21XLTH U12 ( .A0(n7), .A1(n24), .B0(in[6]), .Y(n5) );
  INVXLTH U13 ( .A(in[3]), .Y(n24) );
  XOR2XLTH U14 ( .A(in[0]), .B(n26), .Y(n10) );
  INVXLTH U15 ( .A(in[1]), .Y(n26) );
  OAI221XLTH U17 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n26), .C0(n6), .Y(
        out[1]) );
  OAI221XLTH U18 ( .A0(n29), .A1(n8), .B0(in[6]), .B1(n25), .C0(n6), .Y(out[2]) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  AOI21X8 U5 ( .A0(in[6]), .A1(n11), .B0(n28), .Y(n6) );
  AOI2BB1X4 U16 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n28) );
  INVXLTH U20 ( .A(in[6]), .Y(n29) );
endmodule


module tc_sm_77 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n17, n19, n20, n21, n22, n23, n24,
         n26;

  OAI33X4 U3 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n20), .B2(n21), .Y(n8) );
  INVXLTH U4 ( .A(in[4]), .Y(n21) );
  INVX2TH U5 ( .A(in[5]), .Y(n20) );
  OAI221X2TH U6 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n26), .Y(
        out[1]) );
  OAI33X2 U7 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n20), .B2(n21), .Y(n17) );
  INVXLTH U8 ( .A(in[6]), .Y(n19) );
  OAI221XLTH U9 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2]) );
  OAI2BB1X4 U10 ( .A0N(n22), .A1N(n9), .B0(in[6]), .Y(n13) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n22) );
  XNOR2XLTH U13 ( .A(n23), .B(n11), .Y(n10) );
  OAI21XLTH U14 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n26), .Y(out[0]) );
  INVXLTH U17 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U20 ( .A(in[2]), .Y(n23) );
  OAI211XLTH U21 ( .A0(in[6]), .A1(n22), .B0(n8), .C0(n7), .Y(out[3]) );
  CLKBUFX40 U22 ( .A(n17), .Y(n26) );
endmodule


module tc_sm_76 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n22, n23, n24, n25, n27, n28,
         n29;

  OAI211X1 U3 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221X2TH U4 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[2]) );
  OAI221X1 U5 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[1])
         );
  INVXLTH U6 ( .A(in[6]), .Y(n20) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U10 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U11 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  XNOR2XLTH U12 ( .A(n24), .B(n11), .Y(n10) );
  NAND2BXLTH U13 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVX2 U14 ( .A(in[5]), .Y(n21) );
  INVXLTH U15 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U18 ( .A(in[2]), .Y(n24) );
  INVXL U20 ( .A(in[4]), .Y(n22) );
  AOI33X4 U7 ( .A0(n22), .A1(n28), .A2(n21), .B0(n29), .B1(in[5]), .B2(in[4]), 
        .Y(n27) );
  CLKINVX40 U19 ( .A(n27), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n28) );
  AOI21BX4 U22 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n29) );
endmodule


module total_3_test_28 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n5, n6, n41, n42, n43, n44, n45, n46, n47, n48, n53, n54;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_79 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_78 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_77 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_76 sm_tc_4 ( .out(in1), .in(in) );
  add_19 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_79 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_78 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_77 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_76 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXL up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n44), .CK(clk), .RN(n6), 
        .Q(up1[2]) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n44), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQX1 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n47), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n45), .CK(clk), .RN(n6), .Q(
        h) );
  SDFFRHQX1TH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n42), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  SDFFRHQX1TH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up3[3]) );
  SDFFRHQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n47), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRHQX1TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n44), .CK(clk), .RN(n5), 
        .Q(up3[4]) );
  SDFFRQXLTH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n42), .CK(clk), .RN(n5), 
        .Q(up2[1]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n48), .CK(clk), .RN(n5), .Q(
        up1[0]) );
  SDFFRHQX1TH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n44), .CK(clk), .RN(n5), 
        .Q(up2[2]) );
  SDFFRHQX1TH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n45), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n43), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRHQX2 up3_reg_0_ ( .D(w8[0]), .SI(n54), .SE(n45), .CK(clk), .RN(n5), .Q(
        up3[0]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n6) );
  BUFX3TH U4 ( .A(rst), .Y(n5) );
  SDFFRX4 up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n45), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n43), .CK(clk), .RN(n6), 
        .Q(up1[3]) );
  DLY1X1TH U37 ( .A(n46), .Y(n41) );
  INVXLTH U38 ( .A(n41), .Y(n42) );
  INVXLTH U39 ( .A(n41), .Y(n43) );
  DLY1X1TH U40 ( .A(test_se), .Y(n44) );
  DLY1X1TH U41 ( .A(test_se), .Y(n45) );
  INVXLTH U42 ( .A(test_se), .Y(n46) );
  INVXLTH U43 ( .A(n41), .Y(n47) );
  INVXLTH U44 ( .A(n41), .Y(n48) );
  INVXLTH U45 ( .A(up2[4]), .Y(n53) );
  INVXLTH U46 ( .A(n53), .Y(n54) );
endmodule


module sm_tc_75 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n21, n22, n25, n26;

  XNOR2X2 U2 ( .A(n22), .B(n8), .Y(n5) );
  INVX2 U3 ( .A(in[2]), .Y(n22) );
  AOI31X1 U5 ( .A0(n3), .A1(n4), .A2(n5), .B0(n21), .Y(out[4]) );
  OAI22X1 U6 ( .A0(in[4]), .A1(n22), .B0(n21), .B1(n5), .Y(out[2]) );
  AO21X2 U7 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  BUFX2TH U8 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X4TH U9 ( .B0(n21), .B1(n6), .A0N(in[1]), .A1N(n21), .Y(out[1]) );
  OAI2BB2XLTH U10 ( .B0(n21), .B1(n4), .A0N(in[3]), .A1N(n21), .Y(out[3]) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  INVX3TH U13 ( .A(in[4]), .Y(n21) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  OR2X8 U4 ( .A(in[1]), .B(in[0]), .Y(n25) );
  CLKINVX40 U12 ( .A(n25), .Y(n8) );
  XOR2X1 U14 ( .A(n26), .B(in[3]), .Y(n4) );
  CLKAND2X12 U17 ( .A(n8), .B(n22), .Y(n26) );
endmodule


module sm_tc_74 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n37, n3, n4, n5, n6, n7, n8, n24, n26, n29, n30, n33, n34, n36;

  OAI2BB2X2 U5 ( .B0(n29), .B1(n6), .A0N(in[1]), .A1N(n29), .Y(out[1]) );
  NAND2X2 U2 ( .A(n8), .B(n30), .Y(n7) );
  XNOR2X1TH U3 ( .A(n30), .B(n8), .Y(n5) );
  NOR2BXL U4 ( .AN(n6), .B(n24), .Y(n3) );
  XNOR2X2 U6 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX2TH U7 ( .A(in[4]), .Y(n29) );
  BUFX5 U8 ( .A(in[0]), .Y(n24) );
  INVX2TH U9 ( .A(out[4]), .Y(n26) );
  INVX2 U10 ( .A(in[2]), .Y(n30) );
  AOI31X2TH U11 ( .A0(n3), .A1(n4), .A2(n5), .B0(n29), .Y(n37) );
  OAI22X1 U12 ( .A0(in[4]), .A1(n30), .B0(n29), .B1(n5), .Y(out[2]) );
  AO21XLTH U14 ( .A0(n24), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2XLTH U15 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  INVXLTH U16 ( .A(n26), .Y(out[5]) );
  INVXLTH U17 ( .A(n26), .Y(out[6]) );
  BUFX2TH U18 ( .A(n24), .Y(out[0]) );
  CLKBUFX40 U13 ( .A(n37), .Y(n33) );
  CLKINVX40 U19 ( .A(n33), .Y(n34) );
  CLKINVX40 U20 ( .A(n34), .Y(out[4]) );
  OR2X8 U21 ( .A(in[1]), .B(n24), .Y(n36) );
  CLKINVX40 U22 ( .A(n36), .Y(n8) );
endmodule


module sm_tc_73 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n26, n27, n28, n29, n30, n34, n35, n38, n39, n40;

  INVX2 U2 ( .A(n26), .Y(n34) );
  AO21X1 U3 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  BUFX4 U4 ( .A(in[4]), .Y(n26) );
  BUFX2TH U5 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1 U6 ( .A(n35), .B(n8), .Y(n5) );
  OAI2BB2X2TH U10 ( .B0(n34), .B1(n4), .A0N(in[3]), .A1N(n34), .Y(out[3]) );
  OAI2BB2X2TH U11 ( .B0(n34), .B1(n6), .A0N(in[1]), .A1N(n34), .Y(out[1]) );
  CLKINVX2TH U14 ( .A(n4), .Y(n28) );
  NOR3X4 U15 ( .A(n27), .B(n28), .C(n29), .Y(n30) );
  INVXLTH U16 ( .A(n3), .Y(n27) );
  INVXLTH U17 ( .A(n5), .Y(n29) );
  INVXLTH U19 ( .A(n39), .Y(out[6]) );
  CLKINVX1TH U20 ( .A(in[2]), .Y(n35) );
  NOR2BXLTH U21 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKINVX1TH U22 ( .A(n39), .Y(out[5]) );
  NOR2BX8 U7 ( .AN(n38), .B(out[0]), .Y(n8) );
  CLKINVX40 U8 ( .A(in[1]), .Y(n38) );
  OAI2B2X2 U9 ( .A1N(n26), .A0(n5), .B0(n26), .B1(n35), .Y(out[2]) );
  OR2X8 U12 ( .A(n30), .B(n34), .Y(n39) );
  CLKINVX40 U13 ( .A(n39), .Y(out[4]) );
  XOR2X1 U18 ( .A(n40), .B(in[3]), .Y(n4) );
  CLKAND2X12 U23 ( .A(n8), .B(n35), .Y(n40) );
endmodule


module sm_tc_72 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  AOI31X2 U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  OAI22X1TH U3 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  XNOR2X2TH U4 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX1TH U5 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X2TH U6 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  OAI2BB2XLTH U7 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  NOR2X1TH U8 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U9 ( .A(in[2]), .Y(n21) );
  NAND2XLTH U10 ( .A(n8), .B(n21), .Y(n7) );
  CLKINVX2TH U11 ( .A(in[4]), .Y(n22) );
  INVXLTH U12 ( .A(out[4]), .Y(n18) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U14 ( .A(n18), .Y(out[5]) );
  INVXLTH U15 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U16 ( .A(n21), .B(n8), .Y(n5) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_18_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR2X2TH U1 ( .A(B[6]), .B(A[6]), .Y(n2) );
  CLKXOR2X8 U3 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_18_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n5), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX4TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR2X1 U1 ( .A(n1), .B(A[3]), .Y(SUM[3]) );
  NAND2XL U2 ( .A(A[3]), .B(carry[3]), .Y(n2) );
  NAND2XL U3 ( .A(carry[3]), .B(B[3]), .Y(n4) );
  NAND3X2 U4 ( .A(n2), .B(n3), .C(n4), .Y(carry[4]) );
  NAND2XLTH U5 ( .A(A[3]), .B(B[3]), .Y(n3) );
  XOR2XLTH U6 ( .A(B[3]), .B(carry[3]), .Y(n1) );
  AND2XLTH U7 ( .A(B[0]), .B(A[0]), .Y(n5) );
  CLKXOR2X1TH U8 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_18_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_18_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_18_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX1 U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_18_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2TH U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_18 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35;

  add_18_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in2[6], n30, in2[4], n31, n34, 
        in2[1:0]}), .SUM(out3) );
  add_18_DW01_add_1 add_33 ( .A({temp2_6_, n35, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, n25}), .B({in[6:4], n32, n24, in[1:0]}), .SUM(out1) );
  add_18_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in3[6:3], n27, n33, n26}), .SUM(
        out2) );
  add_18_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({temp2_6_, n35, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, n25}), .SUM(out) );
  add_18_DW01_add_4 add_30 ( .A({in2[6], n29, in2[4], n31, n34, in2[1:0]}), 
        .B({in3[6:3], n27, n33, n26}), .SUM({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_18_DW01_add_5 add_29 ( .A({in[6:4], n32, n24, in[1:0]}), .B(in1), .SUM({
        temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_})
         );
  BUFX2 U1 ( .A(in[2]), .Y(n24) );
  BUFX2TH U2 ( .A(in3[0]), .Y(n26) );
  CLKBUFX1TH U3 ( .A(in3[2]), .Y(n27) );
  BUFX2 U4 ( .A(temp2_0_), .Y(n25) );
  INVX2TH U5 ( .A(in2[5]), .Y(n28) );
  BUFX2TH U6 ( .A(in[3]), .Y(n32) );
  CLKBUFX1TH U13 ( .A(in2[3]), .Y(n31) );
  INVXLTH U14 ( .A(n28), .Y(n29) );
  INVXLTH U15 ( .A(n28), .Y(n30) );
  CLKBUFX40 U16 ( .A(in3[1]), .Y(n33) );
  CLKBUFX40 U17 ( .A(in2[2]), .Y(n34) );
  CLKBUFX40 U18 ( .A(temp2_5_), .Y(n35) );
endmodule


module tc_sm_75 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29, n30;

  CLKBUFX1TH U3 ( .A(in[6]), .Y(out[4]) );
  CLKBUFX2TH U4 ( .A(in[6]), .Y(n24) );
  NOR3X1TH U5 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U6 ( .A(in[1]), .Y(n30) );
  XNOR2XLTH U7 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U8 ( .A(in[2]), .Y(n29) );
  XNOR2XLTH U9 ( .A(n29), .B(n11), .Y(n10) );
  NOR2XLTH U10 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U11 ( .A(n24), .Y(n25) );
  OAI33X4TH U12 ( .A0(in[4]), .A1(n24), .A2(in[5]), .B0(n13), .B1(n26), .B2(
        n27), .Y(n8) );
  INVXLTH U13 ( .A(in[4]), .Y(n27) );
  INVXLTH U14 ( .A(in[5]), .Y(n26) );
  CLKINVX1TH U15 ( .A(in[3]), .Y(n28) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U17 ( .A0(n25), .A1(n12), .B0(n24), .B1(n30), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U18 ( .A0(n25), .A1(n10), .B0(n24), .B1(n29), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U19 ( .A0(n9), .A1(n28), .B0(n24), .Y(n7) );
  OAI211XLTH U20 ( .A0(n24), .A1(n28), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U21 ( .A0N(n28), .A1N(n9), .B0(n24), .Y(n13) );
endmodule


module tc_sm_74 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n21, n22, n23, n25, n26, n27, n28,
         n30, n31;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  DLY2X1TH U3 ( .A(n31), .Y(out[4]) );
  OA21XLTH U4 ( .A0(n31), .A1(n26), .B0(n5), .Y(n21) );
  OAI21XL U6 ( .A0(n7), .A1(n26), .B0(in[6]), .Y(n5) );
  CLKINVX1 U8 ( .A(n31), .Y(n25) );
  INVX2 U9 ( .A(in[3]), .Y(n26) );
  NAND3XL U10 ( .A(n22), .B(n23), .C(n6), .Y(out[2]) );
  XOR2XLTH U11 ( .A(in[2]), .B(n9), .Y(n8) );
  NAND2XLTH U12 ( .A(n21), .B(n6), .Y(out[3]) );
  OR2XLTH U13 ( .A(n25), .B(n8), .Y(n22) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  OAI221XLTH U15 ( .A0(n25), .A1(n10), .B0(n31), .B1(n28), .C0(n6), .Y(out[1])
         );
  OR2XLTH U16 ( .A(n31), .B(n27), .Y(n23) );
  AOI2BB1X4 U17 ( .A0N(in[5]), .A1N(in[4]), .B0(n31), .Y(n12) );
  NOR3X1TH U18 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  INVXLTH U19 ( .A(in[2]), .Y(n27) );
  NOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n9) );
  XOR2XLTH U21 ( .A(in[0]), .B(n28), .Y(n10) );
  INVXLTH U22 ( .A(in[1]), .Y(n28) );
  AO21X4 U5 ( .A0(n31), .A1(n11), .B0(n12), .Y(n30) );
  CLKINVX40 U23 ( .A(n30), .Y(n6) );
  CLKBUFX40 U24 ( .A(in[6]), .Y(n31) );
endmodule


module tc_sm_73 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n18, n19, n20, n22, n23, n24, n25, n26,
         n27;

  CLKINVX6TH U3 ( .A(n18), .Y(n8) );
  NOR3X1TH U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U5 ( .A(in[3]), .Y(n25) );
  INVXLTH U6 ( .A(in[6]), .Y(n22) );
  INVXLTH U7 ( .A(in[5]), .Y(n23) );
  INVXLTH U8 ( .A(in[4]), .Y(n24) );
  AOI21BXLTH U9 ( .A0(n25), .A1(n9), .B0N(in[6]), .Y(n20) );
  INVXLTH U10 ( .A(in[6]), .Y(n19) );
  XNOR2XLTH U11 ( .A(n26), .B(n11), .Y(n10) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI21XLTH U13 ( .A0(n9), .A1(n25), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U15 ( .A(in[1]), .Y(n27) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  AOI33X4 U17 ( .A0(n24), .A1(n19), .A2(n23), .B0(n20), .B1(in[5]), .B2(in[4]), 
        .Y(n18) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U19 ( .A0(n22), .A1(n12), .B0(in[6]), .B1(n27), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U20 ( .A0(n22), .A1(n10), .B0(in[6]), .B1(n26), .C0(n8), .Y(
        out[2]) );
  INVXLTH U21 ( .A(in[2]), .Y(n26) );
  OAI211XLTH U22 ( .A0(in[6]), .A1(n25), .B0(n7), .C0(n8), .Y(out[3]) );
endmodule


module tc_sm_72 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n19, n20, n21, n22, n23, n24;

  INVXLTH U3 ( .A(in[5]), .Y(n20) );
  OAI221X1 U4 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2])
         );
  OAI221X2TH U5 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1]) );
  OAI211X2TH U6 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  CLKINVX1TH U7 ( .A(in[3]), .Y(n22) );
  INVX2TH U8 ( .A(in[4]), .Y(n21) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U10 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n11) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U13 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U14 ( .A(in[1]), .Y(n24) );
  OAI2BB1X4 U15 ( .A0N(n22), .A1N(n9), .B0(in[6]), .Y(n13) );
  INVXLTH U16 ( .A(in[2]), .Y(n23) );
  XNOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U18 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  INVXLTH U19 ( .A(in[6]), .Y(n19) );
  OAI33X4 U20 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n20), .B2(
        n21), .Y(n8) );
endmodule


module total_3_test_29 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n6, n7, n44, n45, n46, n47, n48, n49, n50, n51, n58, n59;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_75 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_74 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_73 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_72 sm_tc_4 ( .out(in1), .in(in) );
  add_18 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_75 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_74 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_73 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_72 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n46), .CK(clk), .RN(n6), 
        .Q(up3[0]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n48), .CK(clk), .RN(n6), .Q(
        up1[0]) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n47), .CK(clk), .RN(n6), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up3[3]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up2[3]) );
  SDFFRHQX4TH up1_reg_4_ ( .D(w6[4]), .SI(n59), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up1[4]) );
  SDFFRQX1TH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up3[1]) );
  SDFFRQX1TH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n45), .CK(clk), .RN(n6), 
        .Q(up2[2]) );
  SDFFRQX1TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n47), .CK(clk), .RN(n6), 
        .Q(up3[4]) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n46), .CK(clk), .RN(n6), 
        .Q(up2[1]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n47), .CK(clk), .RN(n6), 
        .Q(up2[0]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n51), .CK(clk), .RN(n7), 
        .Q(up1[3]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n7) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n6) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up1[2]) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up1[1]) );
  SDFFRX4 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n47), .CK(clk), .RN(n7), 
        .Q(up3[2]) );
  SDFFRX4 h_reg ( .D(w5_4_), .SI(test_si), .SE(n45), .CK(clk), .RN(n7), .Q(h)
         );
  DLY1X1TH U37 ( .A(n49), .Y(n44) );
  INVXLTH U38 ( .A(n44), .Y(n45) );
  INVXLTH U39 ( .A(n44), .Y(n46) );
  DLY1X1TH U40 ( .A(test_se), .Y(n47) );
  DLY1X1TH U41 ( .A(test_se), .Y(n48) );
  INVXLTH U42 ( .A(test_se), .Y(n49) );
  INVXLTH U43 ( .A(n44), .Y(n50) );
  INVXLTH U44 ( .A(n44), .Y(n51) );
  INVXLTH U45 ( .A(up1[3]), .Y(n58) );
  INVXLTH U46 ( .A(n58), .Y(n59) );
endmodule


module sm_tc_71 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n24, n25, n28, n29, n30;

  XNOR2X2 U2 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X4 U3 ( .B0(n29), .B1(n6), .A0N(in[1]), .A1N(n29), .Y(out[1]) );
  NOR2X8 U4 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI22X1 U5 ( .A0(in[4]), .A1(n25), .B0(n29), .B1(n5), .Y(out[2]) );
  OAI2BB2XL U6 ( .B0(n29), .B1(n4), .A0N(in[3]), .A1N(n29), .Y(out[3]) );
  INVX4 U7 ( .A(in[4]), .Y(n24) );
  INVX4 U8 ( .A(in[2]), .Y(n25) );
  AOI31X1 U9 ( .A0(n3), .A1(n4), .A2(n5), .B0(n29), .Y(out[4]) );
  CLKBUFX1TH U11 ( .A(in[0]), .Y(out[0]) );
  AO21X2 U12 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKNAND2X2TH U13 ( .A(n8), .B(n25), .Y(n7) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX40 U10 ( .A(n24), .Y(n28) );
  CLKINVX40 U17 ( .A(n28), .Y(n29) );
  XOR2X1 U18 ( .A(n25), .B(n30), .Y(n5) );
  CLKINVX40 U19 ( .A(n8), .Y(n30) );
endmodule


module sm_tc_70 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n17, n18, n19, n20, n21, n22, n26, n27, n30, n31,
         n32, n33;

  OAI2BB2X1 U2 ( .B0(n27), .B1(n6), .A0N(in[1]), .A1N(n27), .Y(out[1]) );
  BUFX2 U4 ( .A(in[4]), .Y(n18) );
  CLKINVX2 U5 ( .A(n8), .Y(n20) );
  INVX1TH U6 ( .A(in[2]), .Y(n26) );
  AND2XL U7 ( .A(in[0]), .B(in[1]), .Y(n17) );
  AOI31X2TH U9 ( .A0(n3), .A1(n4), .A2(n5), .B0(n27), .Y(out[4]) );
  NAND2X2 U11 ( .A(n21), .B(n22), .Y(n5) );
  CLKNAND2X2TH U12 ( .A(n19), .B(n20), .Y(n22) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[6]) );
  NAND2XL U14 ( .A(n26), .B(n8), .Y(n21) );
  INVXL U15 ( .A(n26), .Y(n19) );
  INVX4 U17 ( .A(n18), .Y(n27) );
  OAI2BB2X1TH U18 ( .B0(n27), .B1(n4), .A0N(in[3]), .A1N(n27), .Y(out[3]) );
  CLKBUFX1TH U20 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U21 ( .AN(n6), .B(in[0]), .Y(n3) );
  BUFX2TH U22 ( .A(in[0]), .Y(out[0]) );
  XOR2X1 U3 ( .A(n30), .B(in[3]), .Y(n4) );
  CLKAND2X12 U8 ( .A(n8), .B(n26), .Y(n30) );
  NAND2BX8 U10 ( .AN(n17), .B(n31), .Y(n6) );
  CLKINVX40 U16 ( .A(n8), .Y(n31) );
  NAND2BX8 U19 ( .AN(in[1]), .B(n33), .Y(n32) );
  CLKINVX40 U23 ( .A(n32), .Y(n8) );
  CLKINVX40 U24 ( .A(in[0]), .Y(n33) );
  AO2B2BX4 U25 ( .A0(n27), .A1N(n26), .B0(n18), .B1N(n5), .Y(out[2]) );
endmodule


module sm_tc_69 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n21, n22, n23, n28, n31;

  NOR2X3TH U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  BUFX2 U4 ( .A(in[4]), .Y(n21) );
  OAI2BB2XL U5 ( .B0(n31), .B1(n4), .A0N(in[3]), .A1N(n31), .Y(out[3]) );
  AOI31X2TH U6 ( .A0(n3), .A1(n4), .A2(n5), .B0(n31), .Y(out[4]) );
  XNOR2X1 U7 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX4 U8 ( .A(in[2]), .Y(n28) );
  CLKNAND2X2TH U10 ( .A(n22), .B(n23), .Y(out[2]) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  OR2XLTH U12 ( .A(n21), .B(n28), .Y(n22) );
  OR2XLTH U13 ( .A(n31), .B(n5), .Y(n23) );
  OAI2BB2X2TH U14 ( .B0(n31), .B1(n6), .A0N(in[1]), .A1N(n31), .Y(out[1]) );
  NAND2XLTH U15 ( .A(n8), .B(n28), .Y(n7) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  AO21XL U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2BXLTH U18 ( .AN(n6), .B(in[0]), .Y(n3) );
  BUFX2TH U19 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1 U3 ( .A(n28), .B(n8), .Y(n5) );
  CLKINVX40 U9 ( .A(n21), .Y(n31) );
endmodule


module sm_tc_68 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  XNOR2X1 U2 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X1TH U3 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U4 ( .A(in[0]), .Y(out[0]) );
  NOR2X4TH U5 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX2TH U6 ( .A(in[4]), .Y(n22) );
  CLKINVX1TH U7 ( .A(in[2]), .Y(n21) );
  AOI31X2TH U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U9 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U10 ( .A(out[4]), .Y(n18) );
  CLKINVX1TH U11 ( .A(n18), .Y(out[5]) );
  OAI22X1TH U12 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  OAI2BB2X1TH U13 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  INVXLTH U14 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U15 ( .A(n21), .B(n8), .Y(n5) );
  NAND2XLTH U16 ( .A(n8), .B(n21), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_17_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_17_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_17_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_17_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_17_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n6, n7, n8, n9;
  wire   [6:2] carry;

  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(carry[3]), .CI(B[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_1 ( .A(B[1]), .B(n1), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  INVXLTH U4 ( .A(B[0]), .Y(n7) );
  INVXLTH U5 ( .A(A[0]), .Y(n6) );
  AND2X8 U1 ( .A(n7), .B(A[0]), .Y(n8) );
  OR2X8 U2 ( .A(n9), .B(n8), .Y(SUM[0]) );
  CLKAND2X12 U6 ( .A(B[0]), .B(n6), .Y(n9) );
endmodule


module add_17_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n2;
  wire   [6:2] carry;

  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR2X3TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n2) );
endmodule


module add_17 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n16, n17, n18, n19;

  add_17_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in2[6:3], n19, n17, in2[0]}), 
        .SUM(out3) );
  add_17_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_17_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in3[6:2], n18, in3[0]}), .SUM(out2) );
  add_17_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, n16, temp2_0_}), .SUM(out) );
  add_17_DW01_add_4 add_30 ( .A({in2[6:3], n19, in2[1:0]}), .B({in3[6:2], n18, 
        in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_17_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2 U1 ( .A(in2[1]), .Y(n17) );
  BUFX2 U2 ( .A(temp2_1_), .Y(n16) );
  CLKBUFX40 U3 ( .A(in3[1]), .Y(n18) );
  CLKBUFX40 U4 ( .A(in2[2]), .Y(n19) );
endmodule


module tc_sm_71 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n28) );
  XNOR2XLTH U7 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXLTH U10 ( .A(in[4]), .Y(n26) );
  INVXLTH U11 ( .A(in[5]), .Y(n25) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n27) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n24) );
  OAI221XLTH U16 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_70 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n20, n21, n22, n23, n24, n25,
         n26;

  OAI221X1 U3 ( .A0(n21), .A1(n12), .B0(in[6]), .B1(n26), .C0(n18), .Y(out[1])
         );
  BUFX10 U4 ( .A(n8), .Y(n18) );
  OAI211XL U5 ( .A0(in[6]), .A1(n24), .B0(n7), .C0(n18), .Y(out[3]) );
  OAI221XL U6 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n25), .C0(n18), .Y(out[2])
         );
  INVXL U7 ( .A(in[6]), .Y(n21) );
  INVXLTH U8 ( .A(in[4]), .Y(n23) );
  INVX2TH U9 ( .A(in[5]), .Y(n22) );
  NAND2BXLTH U10 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  OAI21X8 U11 ( .A0(in[3]), .A1(n20), .B0(in[6]), .Y(n13) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U13 ( .A(n9), .Y(n20) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U15 ( .A(n25), .B(n11), .Y(n10) );
  INVXLTH U16 ( .A(in[2]), .Y(n25) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI21XLTH U18 ( .A0(n9), .A1(n24), .B0(in[6]), .Y(n7) );
  INVXLTH U19 ( .A(in[3]), .Y(n24) );
  INVXLTH U20 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI33X4 U22 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n22), .B2(
        n23), .Y(n8) );
endmodule


module tc_sm_69 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n17, n18, n19, n21, n22, n23, n24, n25;

  CLKINVX8 U3 ( .A(n18), .Y(n8) );
  AOI33X2 U4 ( .A0(n22), .A1(n19), .A2(n21), .B0(n17), .B1(in[5]), .B2(in[4]), 
        .Y(n18) );
  INVX2 U5 ( .A(in[6]), .Y(n19) );
  AOI21BX2TH U6 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n17) );
  INVX2TH U7 ( .A(in[5]), .Y(n21) );
  INVXLTH U8 ( .A(in[4]), .Y(n22) );
  OAI221XLTH U9 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[2]) );
  OAI221XLTH U10 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(
        out[1]) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  OAI21XLTH U13 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  XNOR2XLTH U14 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[2]), .Y(n24) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U18 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211XLTH U21 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
endmodule


module tc_sm_68 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n26, n27,
         n28;

  OAI221X2 U4 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2])
         );
  INVXLTH U5 ( .A(in[6]), .Y(n19) );
  CLKINVX1TH U6 ( .A(in[3]), .Y(n22) );
  NOR3X1TH U7 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U8 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U9 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U10 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U11 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U13 ( .A(in[2]), .Y(n23) );
  OAI21XLTH U14 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  INVX2 U15 ( .A(in[5]), .Y(n20) );
  OAI221XLTH U16 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(
        out[1]) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211XLTH U18 ( .A0(in[6]), .A1(n22), .B0(n8), .C0(n7), .Y(out[3]) );
  INVXL U20 ( .A(in[4]), .Y(n21) );
  AOI33X4 U3 ( .A0(n21), .A1(n27), .A2(n20), .B0(n28), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U19 ( .A(n26), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n27) );
  AOI21BX4 U22 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n28) );
endmodule


module total_3_test_30 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n69, w5_4_, n7, n8, n9, n10, n11, n43, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n67;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_71 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_70 sm_tc_2 ( .out(b1), .in({b[4:1], n9}) );
  sm_tc_69 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_68 sm_tc_4 ( .out(in1), .in(in) );
  add_17 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_71 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_70 tc_sm_2 ( .out(w6), .in({n53, w66[5:0]}) );
  tc_sm_69 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_68 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n61), .CK(clk), .RN(n10), 
        .Q(up2[0]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n56), .CK(clk), .RN(n11), 
        .Q(h) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(n43), .SE(n62), .CK(clk), .RN(n10), 
        .Q(up3[3]) );
  SDFFRQX1TH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n59), .CK(clk), .RN(n10), 
        .Q(up2[2]) );
  SDFFRQX1TH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n57), .CK(clk), .RN(n10), 
        .Q(up3[1]) );
  SDFFRQX2TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n59), .CK(clk), .RN(n10), 
        .Q(up3[4]) );
  SDFFSRXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n57), .CK(clk), .SN(1'b1), .RN(rst), .Q(up3[2]), .QN(n43) );
  SDFFRQXLTH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n58), .CK(clk), .RN(n10), .Q(
        n69) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n62), .CK(clk), .RN(n10), 
        .Q(up1[4]) );
  SDFFRQX2 up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n61), .CK(clk), .RN(n10), 
        .Q(up3[0]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n58), .CK(clk), .RN(n10), 
        .Q(up2[4]) );
  CLKBUFX4 U3 ( .A(b[0]), .Y(n9) );
  BUFX3TH U4 ( .A(rst), .Y(n10) );
  CLKINVX8TH U7 ( .A(n7), .Y(n8) );
  INVX3 U8 ( .A(w66[6]), .Y(n7) );
  CLKBUFX1TH U9 ( .A(rst), .Y(n11) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n59), .CK(clk), .RN(n10), 
        .Q(up1[2]) );
  SDFFRX4 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n58), .CK(clk), .RN(n10), 
        .Q(up2[3]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n59), .CK(clk), .RN(n11), 
        .Q(up1[3]) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n56), .CK(clk), .RN(n11), 
        .Q(up1[1]) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n58), .CK(clk), .RN(n10), 
        .Q(up2[1]) );
  CLKINVX40 U41 ( .A(n8), .Y(n52) );
  CLKINVX40 U42 ( .A(n52), .Y(n53) );
  DLY1X1TH U43 ( .A(n69), .Y(n54) );
  INVXLTH U44 ( .A(test_se), .Y(n55) );
  INVXLTH U45 ( .A(n60), .Y(n56) );
  INVXLTH U46 ( .A(n60), .Y(n57) );
  DLY1X1TH U47 ( .A(test_se), .Y(n58) );
  DLY1X1TH U48 ( .A(test_se), .Y(n59) );
  INVXLTH U49 ( .A(test_se), .Y(n60) );
  INVXLTH U50 ( .A(n55), .Y(n61) );
  INVXLTH U51 ( .A(n55), .Y(n62) );
  CLKINVX40 U52 ( .A(n54), .Y(n67) );
  CLKINVX40 U53 ( .A(n67), .Y(up1[0]) );
endmodule


module sm_tc_67 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n26, n27;

  INVX4 U2 ( .A(in[4]), .Y(n26) );
  CLKBUFX2 U3 ( .A(in[0]), .Y(out[0]) );
  AO21X2 U4 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X6 U5 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X1 U6 ( .A(n27), .B(n8), .Y(n5) );
  NAND2X2 U7 ( .A(n8), .B(n27), .Y(n7) );
  OAI2BB2X4 U8 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n26), .Y(out[1]) );
  CLKBUFX1TH U9 ( .A(out[6]), .Y(out[4]) );
  INVX2TH U10 ( .A(in[2]), .Y(n27) );
  OAI22X2TH U11 ( .A0(in[4]), .A1(n27), .B0(n26), .B1(n5), .Y(out[2]) );
  XNOR2X2TH U12 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2XLTH U13 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U15 ( .A(out[6]), .Y(out[5]) );
  AOI31X2TH U16 ( .A0(n3), .A1(n4), .A2(n5), .B0(n26), .Y(out[6]) );
endmodule


module sm_tc_66 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n20, n21, n24, n25, n26;

  NOR2X2 U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  NAND2XLTH U3 ( .A(n8), .B(n21), .Y(n7) );
  INVX2TH U4 ( .A(in[4]), .Y(n20) );
  OAI2BB2X4TH U5 ( .B0(n20), .B1(n6), .A0N(in[1]), .A1N(n20), .Y(out[1]) );
  INVX2TH U6 ( .A(in[2]), .Y(n21) );
  CLKBUFX2TH U7 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U8 ( .A(out[4]), .Y(out[6]) );
  AO21X2TH U9 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  AOI31X2TH U11 ( .A0(n3), .A1(n4), .A2(n5), .B0(n20), .Y(out[4]) );
  OAI22X2TH U12 ( .A0(in[4]), .A1(n21), .B0(n20), .B1(n5), .Y(out[2]) );
  XNOR2X1TH U13 ( .A(n21), .B(n8), .Y(n5) );
  OAI2BB2X1TH U14 ( .B0(n20), .B1(n4), .A0N(n24), .A1N(n20), .Y(out[3]) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX40 U10 ( .A(in[3]), .Y(n24) );
  DLY1X1TH U17 ( .A(n26), .Y(n25) );
  XOR2X1 U18 ( .A(n7), .B(n24), .Y(n26) );
  CLKINVX40 U19 ( .A(n25), .Y(n4) );
endmodule


module sm_tc_65 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n24, n25, n28, n29, n30, n31;

  OAI2BB2X2 U5 ( .B0(n24), .B1(n6), .A0N(in[1]), .A1N(n24), .Y(out[1]) );
  XNOR2X1 U2 ( .A(n30), .B(n8), .Y(n5) );
  OAI22X1 U3 ( .A0(in[4]), .A1(n30), .B0(n28), .B1(n5), .Y(out[2]) );
  INVX4 U4 ( .A(in[4]), .Y(n24) );
  NOR2X4 U6 ( .A(in[1]), .B(in[0]), .Y(n8) );
  NAND2X1 U9 ( .A(n8), .B(n30), .Y(n7) );
  CLKBUFX1TH U10 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  AOI31X4TH U12 ( .A0(n3), .A1(n4), .A2(n5), .B0(n28), .Y(out[4]) );
  CLKINVX1TH U13 ( .A(in[2]), .Y(n25) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U15 ( .AN(n6), .B(out[0]), .Y(n3) );
  AO21XLTH U16 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKBUFX40 U7 ( .A(n24), .Y(n28) );
  AO2B2X4 U8 ( .B0(in[3]), .B1(n28), .A0(n29), .A1N(n28), .Y(out[3]) );
  DLY1X1TH U17 ( .A(n31), .Y(n29) );
  CLKBUFX40 U18 ( .A(n25), .Y(n30) );
  XOR2X1 U19 ( .A(n7), .B(in[3]), .Y(n31) );
  CLKINVX40 U20 ( .A(n29), .Y(n4) );
endmodule


module sm_tc_64 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n20, n21;

  CLKBUFX1TH U2 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1 U3 ( .A(n20), .B(n8), .Y(n5) );
  NOR2X2TH U4 ( .A(in[1]), .B(in[0]), .Y(n8) );
  AO21X1TH U5 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2X1TH U6 ( .B0(n21), .B1(n4), .A0N(in[3]), .A1N(n21), .Y(out[3]) );
  AOI31X2TH U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n21), .Y(out[6]) );
  XNOR2X2TH U8 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X1TH U9 ( .B0(n21), .B1(n6), .A0N(in[1]), .A1N(n21), .Y(out[1]) );
  NOR2BXLTH U10 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n20) );
  NAND2XLTH U12 ( .A(n8), .B(n20), .Y(n7) );
  CLKINVX2TH U13 ( .A(in[4]), .Y(n21) );
  CLKBUFX1TH U14 ( .A(out[6]), .Y(out[4]) );
  CLKBUFX1TH U15 ( .A(out[6]), .Y(out[5]) );
  OAI22X1TH U16 ( .A0(in[4]), .A1(n20), .B0(n21), .B1(n5), .Y(out[2]) );
endmodule


module add_16_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_16_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3;
  wire   [6:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(carry[3]), .B(B[3]), .CI(A[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  CLKBUFX40 U3 ( .A(n3), .Y(n2) );
  XNOR3X2 U4 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n3) );
  CLKINVX40 U5 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_16_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_16_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_16_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_16_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n2;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(B[1]), .B(n2), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n2) );
  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_16 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n25, n26, n27, n28, n29, n30, n31;

  add_16_DW01_add_0 add_34 ( .A({temp1_6_, n30, temp1_4_, n31, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in2[6:4], n29, in2[2:0]}), .SUM(out3) );
  add_16_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, n28, temp2_0_}), .B(in), .SUM(out1) );
  add_16_DW01_add_2 add_32 ( .A({temp1_6_, n30, temp1_4_, n31, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in3[6:3], n27, in3[1], n26}), .SUM(out2) );
  add_16_DW01_add_3 add_31 ( .A({temp1_6_, n30, temp1_4_, n31, temp1_2_, 
        temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, n28, temp2_0_}), .SUM(out) );
  add_16_DW01_add_4 add_30 ( .A({in2[6:4], n29, in2[2:0]}), .B({in3[6:3], n27, 
        in3[1:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_16_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  INVXLTH U1 ( .A(in3[0]), .Y(n25) );
  INVXLTH U2 ( .A(n25), .Y(n26) );
  BUFX3 U3 ( .A(in3[2]), .Y(n27) );
  CLKBUFX40 U4 ( .A(temp2_1_), .Y(n28) );
  CLKBUFX40 U5 ( .A(in2[3]), .Y(n29) );
  CLKBUFX40 U6 ( .A(temp1_5_), .Y(n30) );
  CLKBUFX40 U13 ( .A(temp1_3_), .Y(n31) );
endmodule


module tc_sm_67 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(in[6]), .Y(n26) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n28) );
  INVXLTH U12 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI2BB1XLTH U19 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI211XLTH U20 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
endmodule


module tc_sm_66 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n31, n35, n36, n37, n38, n40, n41,
         n42;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[5]), .C0(in[4]), .Y(n11) );
  OAI221XL U3 ( .A0(n35), .A1(n8), .B0(in[6]), .B1(n37), .C0(n6), .Y(out[2])
         );
  CLKINVX1 U4 ( .A(in[6]), .Y(n35) );
  NOR2X4TH U6 ( .A(n35), .B(n10), .Y(n31) );
  AOI21X8 U8 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n6) );
  XOR2XLTH U10 ( .A(in[0]), .B(n38), .Y(n10) );
  AOI2BB1X4 U13 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  NOR3X1TH U15 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U16 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  INVXLTH U18 ( .A(in[3]), .Y(n36) );
  INVXLTH U19 ( .A(in[1]), .Y(n38) );
  INVXLTH U20 ( .A(in[2]), .Y(n37) );
  XOR2XLTH U21 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U22 ( .A(in[0]), .B(in[1]), .Y(n9) );
  NAND3BX4 U5 ( .AN(n31), .B(n40), .C(n6), .Y(out[1]) );
  OR2X8 U9 ( .A(in[6]), .B(n38), .Y(n40) );
  OAI2B11X4 U11 ( .A1N(n41), .A0(n36), .B0(n5), .C0(n6), .Y(out[3]) );
  CLKINVX40 U12 ( .A(in[6]), .Y(n41) );
  OA21X4 U14 ( .A0(n7), .A1(n36), .B0(in[6]), .Y(n42) );
  CLKINVX40 U23 ( .A(n42), .Y(n5) );
endmodule


module tc_sm_65 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n23, n24, n25, n27, n28, n29,
         n30, n31, n32;

  OAI211X1TH U5 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221XL U6 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[1])
         );
  OAI221XL U7 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[2])
         );
  INVX2TH U8 ( .A(in[5]), .Y(n21) );
  INVXLTH U9 ( .A(in[6]), .Y(n20) );
  CLKINVX1TH U10 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U12 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U14 ( .A(in[2]), .Y(n24) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U16 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U18 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  DLY1X1TH U3 ( .A(in[4]), .Y(n27) );
  AOI33X4 U4 ( .A0(n29), .A1(n30), .A2(n21), .B0(n32), .B1(n31), .B2(in[4]), 
        .Y(n28) );
  CLKINVX40 U20 ( .A(n28), .Y(n8) );
  CLKINVX40 U21 ( .A(n27), .Y(n29) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n30) );
  CLKINVX40 U23 ( .A(n21), .Y(n31) );
  AOI21BX4 U24 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n32) );
endmodule


module tc_sm_64 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n21, n22, n24, n25, n26, n28, n29, n30,
         n31, n32;

  OAI211XLTH U6 ( .A0(in[6]), .A1(n24), .B0(n7), .C0(n8), .Y(out[3]) );
  CLKINVX1TH U7 ( .A(in[3]), .Y(n24) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U9 ( .A(n25), .B(n11), .Y(n10) );
  INVXLTH U10 ( .A(in[2]), .Y(n25) );
  NOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U12 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U14 ( .A0(n9), .A1(n24), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  INVX2 U16 ( .A(in[5]), .Y(n22) );
  OAI221XLTH U17 ( .A0(n21), .A1(n12), .B0(in[6]), .B1(n26), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U18 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n25), .C0(n8), .Y(
        out[2]) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U20 ( .A(in[6]), .Y(n21) );
  INVXLTH U3 ( .A(n30), .Y(n28) );
  AOI33X4 U4 ( .A0(n30), .A1(n31), .A2(n22), .B0(n32), .B1(in[5]), .B2(n28), 
        .Y(n29) );
  CLKINVX40 U5 ( .A(n29), .Y(n8) );
  CLKINVX40 U21 ( .A(in[4]), .Y(n30) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n31) );
  AOI21BX4 U23 ( .A0(n24), .A1(n9), .B0N(in[6]), .Y(n32) );
endmodule


module total_3_test_31 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n6, n7, n44, n45, n46, n47, n48, n49, n50, n51;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_67 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_66 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_65 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_64 sm_tc_4 ( .out(in1), .in(in) );
  add_16 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_67 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_66 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_65 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_64 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n46), .CK(clk), .RN(n6), 
        .Q(up3[3]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up3[0]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up1[3]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n50), .CK(clk), .RN(n7), .Q(
        h) );
  SDFFRHQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n48), .CK(clk), .RN(n7), 
        .Q(up1[4]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n45), .CK(clk), .RN(n6), 
        .Q(up2[4]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n47), .CK(clk), .RN(n6), 
        .Q(up2[3]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n46), .CK(clk), .RN(n6), 
        .Q(up2[0]) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up2[1]) );
  SDFFRQX1TH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n47), .CK(clk), .RN(n6), 
        .Q(up2[2]) );
  SDFFRQX2 up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n47), .CK(clk), .RN(n7), 
        .Q(up3[4]) );
  SDFFRQX2 up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n48), .CK(clk), .RN(n6), .Q(
        up1[0]) );
  CLKBUFX4TH U3 ( .A(rst), .Y(n6) );
  CLKBUFX1TH U4 ( .A(rst), .Y(n7) );
  SDFFRX4 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n51), .CK(clk), .RN(n6), 
        .Q(up3[2]) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up1[1]) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n47), .CK(clk), .RN(n6), 
        .Q(up3[1]) );
  SDFFRHQX8 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n45), .CK(clk), .RN(n6), 
        .Q(up1[2]) );
  DLY1X1TH U37 ( .A(n49), .Y(n44) );
  INVXLTH U38 ( .A(n44), .Y(n45) );
  INVXLTH U39 ( .A(n44), .Y(n46) );
  DLY1X1TH U40 ( .A(test_se), .Y(n47) );
  DLY1X1TH U41 ( .A(test_se), .Y(n48) );
  INVXLTH U42 ( .A(test_se), .Y(n49) );
  INVXLTH U43 ( .A(n44), .Y(n50) );
  INVXLTH U44 ( .A(n44), .Y(n51) );
endmodule


module sm_tc_63 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n22, n23, n24, n25, n26, n30, n31, n34, n35, n36,
         n37, n38, n39;

  AO21X2 U2 ( .A0(in[0]), .A1(n39), .B0(n8), .Y(n6) );
  BUFX2 U3 ( .A(in[0]), .Y(out[0]) );
  AND3X2 U5 ( .A(n3), .B(n4), .C(n5), .Y(n22) );
  NOR2X3 U6 ( .A(n22), .B(n37), .Y(out[4]) );
  INVX6 U8 ( .A(in[4]), .Y(n30) );
  NAND2X2 U9 ( .A(n25), .B(n26), .Y(n5) );
  NAND2X4 U11 ( .A(n23), .B(n24), .Y(n26) );
  CLKINVX1 U12 ( .A(n31), .Y(n23) );
  INVXLTH U13 ( .A(n8), .Y(n24) );
  INVX2 U14 ( .A(in[2]), .Y(n31) );
  OAI22XL U15 ( .A0(n36), .A1(n31), .B0(n37), .B1(n5), .Y(out[2]) );
  OAI2BB2X4 U16 ( .B0(n37), .B1(n6), .A0N(n39), .A1N(n37), .Y(out[1]) );
  CLKBUFX1TH U18 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2XLTH U19 ( .B0(n37), .B1(n4), .A0N(in[3]), .A1N(n37), .Y(out[3]) );
  CLKBUFX1TH U20 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U21 ( .AN(n6), .B(in[0]), .Y(n3) );
  NOR2BX8 U4 ( .AN(n34), .B(in[0]), .Y(n8) );
  CLKINVX40 U7 ( .A(n39), .Y(n34) );
  AND2X8 U10 ( .A(n31), .B(n8), .Y(n35) );
  CLKINVX40 U17 ( .A(n35), .Y(n25) );
  CLKINVX40 U22 ( .A(n30), .Y(n36) );
  CLKINVX40 U23 ( .A(n36), .Y(n37) );
  XOR2X1 U24 ( .A(n38), .B(in[3]), .Y(n4) );
  CLKAND2X12 U25 ( .A(n8), .B(n31), .Y(n38) );
  CLKBUFX40 U26 ( .A(in[1]), .Y(n39) );
endmodule


module sm_tc_62 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n33, n3, n4, n5, n6, n8, n20, n22, n25, n26, n29, n30, n31;

  NOR2X2 U2 ( .A(n31), .B(in[0]), .Y(n8) );
  NOR2BXLTH U3 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX8 U5 ( .A(n20), .Y(n25) );
  CLKBUFX1TH U6 ( .A(in[4]), .Y(n20) );
  CLKBUFX1TH U7 ( .A(in[0]), .Y(out[0]) );
  AOI31X1 U8 ( .A0(n5), .A1(n4), .A2(n3), .B0(n25), .Y(n33) );
  OAI22X1 U9 ( .A0(n20), .A1(n26), .B0(n25), .B1(n5), .Y(out[2]) );
  INVX2 U10 ( .A(in[2]), .Y(n26) );
  INVX2TH U11 ( .A(n33), .Y(n22) );
  AO21XLTH U13 ( .A0(in[0]), .A1(n31), .B0(n8), .Y(n6) );
  OAI2BB2X1TH U14 ( .B0(n25), .B1(n4), .A0N(in[3]), .A1N(n25), .Y(out[3]) );
  INVXLTH U15 ( .A(n22), .Y(out[5]) );
  INVXLTH U16 ( .A(n22), .Y(out[6]) );
  XNOR2X1 U4 ( .A(n26), .B(n8), .Y(n5) );
  XOR2X1 U12 ( .A(n29), .B(in[3]), .Y(n4) );
  CLKAND2X12 U17 ( .A(n8), .B(n26), .Y(n29) );
  AO2B2X4 U18 ( .B0(n31), .B1(n25), .A0(n30), .A1N(n6), .Y(out[1]) );
  CLKINVX40 U19 ( .A(n25), .Y(n30) );
  CLKBUFX40 U20 ( .A(in[1]), .Y(n31) );
  CLKINVX40 U21 ( .A(n22), .Y(out[4]) );
endmodule


module sm_tc_61 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n30, n3, n4, n5, n6, n7, n8, n19, n20, n24, n25, n28;

  NOR2XLTH U2 ( .A(in[4]), .B(n25), .Y(n19) );
  NOR2X1 U3 ( .A(n24), .B(n5), .Y(n20) );
  OR2X2 U4 ( .A(n19), .B(n20), .Y(out[2]) );
  INVX4 U5 ( .A(in[4]), .Y(n24) );
  XNOR2X1 U6 ( .A(n25), .B(n8), .Y(n5) );
  OAI2BB2XL U7 ( .B0(n24), .B1(n4), .A0N(in[3]), .A1N(n24), .Y(out[3]) );
  NAND2X2 U8 ( .A(n8), .B(n25), .Y(n7) );
  NOR2X4 U9 ( .A(in[1]), .B(in[0]), .Y(n8) );
  BUFX2TH U10 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1TH U11 ( .A(n7), .B(in[3]), .Y(n4) );
  AO21X1 U12 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2X2 U13 ( .B0(n24), .B1(n6), .A0N(in[1]), .A1N(n24), .Y(out[1]) );
  INVX1TH U14 ( .A(in[2]), .Y(n25) );
  DLY2X1TH U15 ( .A(out[4]), .Y(out[5]) );
  DLY2X1TH U16 ( .A(out[4]), .Y(out[6]) );
  AOI31X2TH U17 ( .A0(n3), .A1(n4), .A2(n5), .B0(n24), .Y(n30) );
  NOR2BXLTH U18 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKINVX40 U19 ( .A(n30), .Y(n28) );
  CLKINVX40 U20 ( .A(n28), .Y(out[4]) );
endmodule


module sm_tc_60 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22, n25;

  XNOR2X1 U2 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X1TH U3 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  INVXLTH U4 ( .A(n18), .Y(out[5]) );
  OAI22X1TH U5 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  CLKBUFX1TH U6 ( .A(in[0]), .Y(out[0]) );
  NAND2X1TH U7 ( .A(n8), .B(n21), .Y(n7) );
  CLKINVX2TH U8 ( .A(in[4]), .Y(n22) );
  CLKINVX1TH U10 ( .A(in[2]), .Y(n21) );
  INVXLTH U11 ( .A(out[4]), .Y(n18) );
  AOI31X2TH U12 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2BB2X1TH U14 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  INVXLTH U15 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U16 ( .A(n21), .B(n8), .Y(n5) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OR2X8 U9 ( .A(in[1]), .B(in[0]), .Y(n25) );
  CLKINVX40 U18 ( .A(n25), .Y(n8) );
endmodule


module add_15_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR2X1TH U1 ( .A(B[6]), .B(A[6]), .Y(n2) );
  CLKAND2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  CLKXOR2X8 U4 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
endmodule


module add_15_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  ADDFHX2TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKNAND2X2TH U1 ( .A(A[1]), .B(B[1]), .Y(n4) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND3X2TH U3 ( .A(n3), .B(n4), .C(n5), .Y(carry[2]) );
  CLKNAND2X2 U4 ( .A(n1), .B(B[1]), .Y(n5) );
  CLKNAND2X2 U5 ( .A(A[1]), .B(n1), .Y(n3) );
  CLKXOR2X1TH U6 ( .A(n2), .B(A[1]), .Y(SUM[1]) );
  XOR2XLTH U7 ( .A(B[1]), .B(n1), .Y(n2) );
  AND2X1TH U8 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_15_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_15_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_15_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_15_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X4TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_15 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n20, n21, n22, n23, n24, n25, n26, n27, n28;

  add_15_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n25, n28, 
        temp1_1_, temp1_0_}), .B({in2[6:2], n27, in2[0]}), .SUM(out3) );
  add_15_DW01_add_1 add_33 ( .A({temp2_6_, n26, temp2_4_, n21, temp2_2_, 
        temp2_1_, temp2_0_}), .B({in[6:2], n20, in[0]}), .SUM(out1) );
  add_15_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n25, n28, 
        temp1_1_, temp1_0_}), .B({in3[6:4], n24, n23, in3[1:0]}), .SUM(out2)
         );
  add_15_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n25, n28, 
        temp1_1_, temp1_0_}), .B({temp2_6_, n26, temp2_4_, n21, temp2_2_, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_15_DW01_add_4 add_30 ( .A({in2[6:2], n27, in2[0]}), .B({in3[6:4], n24, 
        n23, in3[1:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}) );
  add_15_DW01_add_5 add_29 ( .A({in[6:2], n20, in[0]}), .B(in1), .SUM({
        temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_})
         );
  BUFX2 U1 ( .A(in[1]), .Y(n20) );
  INVX2 U2 ( .A(in3[2]), .Y(n22) );
  INVX2 U3 ( .A(n22), .Y(n23) );
  CLKBUFX2TH U4 ( .A(temp2_3_), .Y(n21) );
  CLKBUFX40 U5 ( .A(in3[3]), .Y(n24) );
  CLKBUFX40 U6 ( .A(temp1_3_), .Y(n25) );
  CLKBUFX40 U13 ( .A(temp2_5_), .Y(n26) );
  CLKBUFX40 U14 ( .A(in2[1]), .Y(n27) );
  CLKBUFX40 U15 ( .A(temp1_2_), .Y(n28) );
endmodule


module tc_sm_63 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n25, n27, n28, n29, n30, n31, n32;

  CLKBUFX2TH U3 ( .A(in[6]), .Y(n25) );
  NOR3X1TH U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U5 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U6 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U7 ( .A(in[2]), .Y(n31) );
  XNOR2XLTH U8 ( .A(n31), .B(n11), .Y(n10) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U10 ( .A(n25), .Y(n27) );
  OAI33X4TH U11 ( .A0(in[4]), .A1(n25), .A2(in[5]), .B0(n13), .B1(n28), .B2(
        n29), .Y(n8) );
  INVXLTH U12 ( .A(in[4]), .Y(n29) );
  INVXLTH U13 ( .A(in[5]), .Y(n28) );
  CLKINVX1TH U14 ( .A(in[3]), .Y(n30) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U17 ( .A0(n27), .A1(n12), .B0(n25), .B1(n32), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U18 ( .A0(n27), .A1(n10), .B0(n25), .B1(n31), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U19 ( .A0(n9), .A1(n30), .B0(n25), .Y(n7) );
  OAI211XLTH U20 ( .A0(n25), .A1(n30), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U21 ( .A0N(n30), .A1N(n9), .B0(n25), .Y(n13) );
endmodule


module tc_sm_62 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n19, n20, n21, n23, n24, n25, n26, n27,
         n28, n30;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  CLKINVX2 U4 ( .A(in[6]), .Y(n25) );
  NAND3XL U5 ( .A(n19), .B(n20), .C(n6), .Y(out[1]) );
  OR2XL U6 ( .A(n25), .B(n10), .Y(n19) );
  AOI21BX4 U8 ( .A0(in[6]), .A1(n11), .B0N(n21), .Y(n6) );
  OAI211X2TH U9 ( .A0(in[6]), .A1(n26), .B0(n5), .C0(n6), .Y(out[3]) );
  NAND3XL U10 ( .A(n23), .B(n24), .C(n6), .Y(out[2]) );
  XOR2XLTH U11 ( .A(in[0]), .B(n28), .Y(n10) );
  OR2XLTH U12 ( .A(in[6]), .B(n28), .Y(n20) );
  OR2X2 U13 ( .A(n25), .B(n8), .Y(n23) );
  XOR2XLTH U14 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR3X1TH U15 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  OAI21XLTH U16 ( .A0(n7), .A1(n26), .B0(in[6]), .Y(n5) );
  INVXLTH U17 ( .A(in[3]), .Y(n26) );
  CLKBUFX1TH U18 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U19 ( .A(in[1]), .Y(n28) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  INVXLTH U21 ( .A(in[2]), .Y(n27) );
  NOR2XLTH U22 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OR2XLTH U23 ( .A(in[6]), .B(n27), .Y(n24) );
  AOI2BB1X4 U3 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n30) );
  CLKINVX40 U24 ( .A(n30), .Y(n21) );
endmodule


module tc_sm_61 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n18, n19, n20, n22, n23, n24, n25, n26,
         n28, n29;

  AOI33X2 U3 ( .A0(n23), .A1(n29), .A2(n22), .B0(n20), .B1(in[5]), .B2(in[4]), 
        .Y(n18) );
  CLKINVX4 U4 ( .A(n18), .Y(n8) );
  OAI221X1 U5 ( .A0(n29), .A1(n10), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[2])
         );
  INVXLTH U6 ( .A(in[5]), .Y(n22) );
  CLKINVX1 U7 ( .A(in[6]), .Y(n19) );
  AOI21BXLTH U8 ( .A0(n24), .A1(n9), .B0N(in[6]), .Y(n20) );
  INVXLTH U9 ( .A(in[4]), .Y(n23) );
  CLKINVX1TH U10 ( .A(in[3]), .Y(n24) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U13 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U15 ( .A(n25), .B(n11), .Y(n10) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U17 ( .A(in[2]), .Y(n25) );
  OAI21XLTH U18 ( .A0(n9), .A1(n24), .B0(in[6]), .Y(n7) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U20 ( .A0(n29), .A1(n12), .B0(in[6]), .B1(n26), .C0(n8), .Y(
        out[1]) );
  CLKINVX40 U21 ( .A(n19), .Y(n28) );
  CLKINVX40 U22 ( .A(n28), .Y(n29) );
  OAI2B11X4 U23 ( .A1N(n29), .A0(n24), .B0(n7), .C0(n8), .Y(out[3]) );
endmodule


module tc_sm_60 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n18, n19, n20, n21, n22, n23, n25, n26,
         n27;

  OAI221XL U3 ( .A0(n18), .A1(n10), .B0(in[6]), .B1(n22), .C0(n8), .Y(out[2])
         );
  OAI221XL U4 ( .A0(n18), .A1(n12), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[1])
         );
  INVXLTH U5 ( .A(in[4]), .Y(n20) );
  INVXLTH U6 ( .A(in[5]), .Y(n19) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n21) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U10 ( .A(in[1]), .Y(n23) );
  XNOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U12 ( .A(n22), .B(n11), .Y(n10) );
  NOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U14 ( .A(in[2]), .Y(n22) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211XLTH U17 ( .A0(in[6]), .A1(n21), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n21), .B0(in[6]), .Y(n7) );
  INVXLTH U19 ( .A(in[6]), .Y(n18) );
  AOI33X4 U7 ( .A0(n20), .A1(n26), .A2(n19), .B0(n27), .B1(in[5]), .B2(in[4]), 
        .Y(n25) );
  CLKINVX40 U20 ( .A(n25), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n26) );
  AOI21BX4 U22 ( .A0(n21), .A1(n9), .B0N(in[6]), .Y(n27) );
endmodule


module total_3_test_32 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n4, n5, n6, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_63 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_62 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_61 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_60 sm_tc_4 ( .out(in1), .in(in) );
  add_15 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_63 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_62 tc_sm_2 ( .out(w6), .in({n4, w66[5:0]}) );
  tc_sm_61 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_60 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up3[3]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n55), .CK(clk), .RN(n5), 
        .Q(up1[3]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n54), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n47), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRQX2TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up3[4]) );
  SDFFRQX1TH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up2[2]) );
  SDFFRQXL up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n55), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n47), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQX2 up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n53), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  BUFX20 U3 ( .A(w66[6]), .Y(n4) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n5) );
  CLKBUFX1TH U5 ( .A(rst), .Y(n6) );
  SDFFRX4 h_reg ( .D(w5_4_), .SI(test_si), .SE(n53), .CK(clk), .RN(n6), .Q(h)
         );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n47), .CK(clk), .RN(n6), 
        .Q(up1[2]) );
  SDFFRHQX8 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up2[1]) );
  SDFFRX4 up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n54), .CK(clk), .RN(n6), .Q(
        up1[0]) );
  DLY1X1TH U38 ( .A(n49), .Y(n46) );
  DLY1X1TH U39 ( .A(n50), .Y(n47) );
  DLY1X1TH U40 ( .A(n52), .Y(n48) );
  INVXLTH U41 ( .A(n48), .Y(n49) );
  INVXLTH U42 ( .A(n52), .Y(n50) );
  DLY1X1TH U43 ( .A(test_se), .Y(n51) );
  INVXLTH U44 ( .A(test_se), .Y(n52) );
  INVXLTH U45 ( .A(n48), .Y(n53) );
  INVXLTH U46 ( .A(n48), .Y(n54) );
  INVXLTH U47 ( .A(n48), .Y(n55) );
endmodule


module sm_tc_59 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n21, n22, n25, n26;

  OAI22XL U2 ( .A0(in[4]), .A1(n22), .B0(n21), .B1(n5), .Y(out[2]) );
  AOI31X1 U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n21), .Y(out[4]) );
  XNOR2X1 U4 ( .A(n7), .B(n26), .Y(n4) );
  AO21XL U5 ( .A0(n25), .A1(in[1]), .B0(n8), .Y(n6) );
  NAND2XLTH U6 ( .A(n8), .B(n22), .Y(n7) );
  OAI2BB2X4 U7 ( .B0(n21), .B1(n6), .A0N(in[1]), .A1N(n21), .Y(out[1]) );
  INVX2TH U8 ( .A(in[2]), .Y(n22) );
  INVX4TH U9 ( .A(in[4]), .Y(n21) );
  CLKBUFX1TH U10 ( .A(n25), .Y(out[0]) );
  OAI2BB2X2TH U11 ( .B0(n21), .B1(n4), .A0N(n26), .A1N(n21), .Y(out[3]) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[5]) );
  NOR2X6 U14 ( .A(in[1]), .B(n25), .Y(n8) );
  NOR2BXLTH U15 ( .AN(n6), .B(n25), .Y(n3) );
  XNOR2X1 U16 ( .A(n22), .B(n8), .Y(n5) );
  CLKBUFX40 U17 ( .A(in[0]), .Y(n25) );
  CLKBUFX40 U18 ( .A(in[3]), .Y(n26) );
endmodule


module sm_tc_58 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n19, n22, n23;

  INVX2 U2 ( .A(in[2]), .Y(n23) );
  XNOR2X1TH U3 ( .A(n7), .B(in[3]), .Y(n4) );
  AOI31X2 U4 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  OAI2BB2XL U5 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  OAI2BB2X2 U6 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  NOR2X2 U7 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX3 U8 ( .A(in[4]), .Y(n22) );
  OAI22X4TH U9 ( .A0(in[4]), .A1(n23), .B0(n22), .B1(n5), .Y(out[2]) );
  INVXLTH U10 ( .A(n19), .Y(out[6]) );
  INVXLTH U11 ( .A(out[4]), .Y(n19) );
  INVXLTH U12 ( .A(n19), .Y(out[5]) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  XNOR2X1TH U14 ( .A(n23), .B(n8), .Y(n5) );
  BUFX2TH U15 ( .A(in[0]), .Y(out[0]) );
  NAND2XLTH U16 ( .A(n8), .B(n23), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module sm_tc_57 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n30, n32, n33, n35, n36, n37;

  AOI31X4 U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n32), .Y(out[6]) );
  CLKBUFX1TH U3 ( .A(out[6]), .Y(out[4]) );
  BUFX2TH U4 ( .A(out[6]), .Y(out[5]) );
  CLKINVX6TH U5 ( .A(n30), .Y(out[0]) );
  INVX1TH U6 ( .A(in[0]), .Y(n30) );
  XNOR2X4 U8 ( .A(n7), .B(in[3]), .Y(n4) );
  NOR2X6TH U9 ( .A(in[1]), .B(out[0]), .Y(n8) );
  AO21X1TH U11 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKINVX1TH U12 ( .A(in[2]), .Y(n33) );
  INVX2TH U13 ( .A(in[4]), .Y(n32) );
  NOR2BXLTH U14 ( .AN(n6), .B(out[0]), .Y(n3) );
  OAI2BB2X1TH U15 ( .B0(n32), .B1(n4), .A0N(in[3]), .A1N(n32), .Y(out[3]) );
  OAI22X4 U16 ( .A0(in[4]), .A1(n37), .B0(n32), .B1(n5), .Y(out[2]) );
  OAI2BB2X4 U17 ( .B0(n32), .B1(n6), .A0N(in[1]), .A1N(n32), .Y(out[1]) );
  XOR2X1 U7 ( .A(n36), .B(n8), .Y(n5) );
  AND2X8 U10 ( .A(n8), .B(n37), .Y(n35) );
  CLKINVX40 U18 ( .A(n35), .Y(n7) );
  CLKINVX40 U19 ( .A(n33), .Y(n36) );
  CLKINVX40 U20 ( .A(n36), .Y(n37) );
endmodule


module sm_tc_56 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n18, n19, n20, n22, n25, n26;

  CLKNAND2X2 U2 ( .A(n7), .B(in[3]), .Y(n19) );
  NAND2X4 U3 ( .A(n17), .B(n18), .Y(n20) );
  NAND2X6 U4 ( .A(n19), .B(n20), .Y(n4) );
  CLKINVX2 U5 ( .A(n7), .Y(n17) );
  INVX2 U6 ( .A(in[3]), .Y(n18) );
  OAI2BB2X4 U7 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  AOI31X2 U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n26), .Y(out[4]) );
  OAI22X2TH U9 ( .A0(in[4]), .A1(n25), .B0(n26), .B1(n5), .Y(out[2]) );
  CLKBUFX1TH U10 ( .A(in[0]), .Y(out[0]) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n25) );
  INVXLTH U12 ( .A(out[4]), .Y(n22) );
  OAI2BB2X1TH U13 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n26), .Y(out[1]) );
  INVXLTH U14 ( .A(n22), .Y(out[6]) );
  NOR2X3TH U15 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX2TH U16 ( .A(in[4]), .Y(n26) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX2TH U18 ( .A(n22), .Y(out[5]) );
  XNOR2X1TH U19 ( .A(n25), .B(n8), .Y(n5) );
  NAND2XLTH U20 ( .A(n8), .B(n25), .Y(n7) );
  AO21XLTH U21 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_14_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_14_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22;
  wire   [5:2] carry;

  ADDFHX4TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  NAND2X2TH U2 ( .A(B[5]), .B(n16), .Y(n4) );
  NAND2XLTH U3 ( .A(A[5]), .B(B[5]), .Y(n13) );
  NAND2XLTH U4 ( .A(carry[5]), .B(A[5]), .Y(n11) );
  INVX2 U6 ( .A(A[5]), .Y(n16) );
  CLKXOR2X4 U8 ( .A(n10), .B(carry[5]), .Y(SUM[5]) );
  CLKNAND2X4TH U9 ( .A(n9), .B(n14), .Y(carry[4]) );
  XOR2X1TH U10 ( .A(B[3]), .B(carry[3]), .Y(n6) );
  NAND2X3TH U11 ( .A(A[3]), .B(carry[3]), .Y(n7) );
  NAND2X4TH U12 ( .A(A[3]), .B(B[3]), .Y(n8) );
  CLKXOR2X1TH U13 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U14 ( .A(B[0]), .B(A[0]), .Y(n1) );
  NAND2XLTH U15 ( .A(carry[5]), .B(B[5]), .Y(n12) );
  XOR2X1TH U17 ( .A(n6), .B(A[3]), .Y(SUM[3]) );
  AND3X2 U19 ( .A(n11), .B(n12), .C(n13), .Y(n15) );
  INVXL U20 ( .A(B[5]), .Y(n17) );
  AND2X8 U1 ( .A(carry[3]), .B(B[3]), .Y(n18) );
  CLKINVX40 U5 ( .A(n18), .Y(n9) );
  AND2X8 U7 ( .A(n17), .B(A[5]), .Y(n19) );
  CLKINVX40 U16 ( .A(n19), .Y(n5) );
  AND2X8 U18 ( .A(n4), .B(n5), .Y(n20) );
  CLKINVX40 U21 ( .A(n20), .Y(n10) );
  NAND2X8 U22 ( .A(n8), .B(n7), .Y(n21) );
  CLKINVX40 U23 ( .A(n21), .Y(n14) );
  XOR3X2 U24 ( .A(A[6]), .B(B[6]), .C(n15), .Y(n22) );
  CLKINVX40 U25 ( .A(n22), .Y(SUM[6]) );
endmodule


module add_14_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2XL U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_14_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(n2), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKINVX40 U4 ( .A(A[6]), .Y(n2) );
endmodule


module add_14_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n7, n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  ADDFX4TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(n7) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  NAND3X4 U1 ( .A(n2), .B(n3), .C(n4), .Y(carry[3]) );
  CLKNAND2X2TH U2 ( .A(carry[2]), .B(B[2]), .Y(n3) );
  CLKNAND2X4 U3 ( .A(carry[2]), .B(A[2]), .Y(n2) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U5 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2XL U6 ( .A(A[2]), .B(B[2]), .Y(n4) );
  XOR3X4TH U7 ( .A(carry[2]), .B(A[2]), .C(B[2]), .Y(SUM[2]) );
  CLKINVX40 U8 ( .A(n7), .Y(n5) );
  CLKINVX40 U9 ( .A(n5), .Y(SUM[5]) );
endmodule


module add_14_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n2;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2TH U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n2) );
endmodule


module add_14 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n19, n20, n21, n22, n23, n24;

  add_14_DW01_add_0 add_34 ( .A({temp1_6_, n24, temp1_4_, temp1_3_, temp1_2_, 
        temp1_1_, n22}), .B({in2[6:4], n23, in2[2], n19, in2[0]}), .SUM(out3)
         );
  add_14_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_14_DW01_add_2 add_32 ( .A({temp1_6_, n24, temp1_4_, temp1_3_, temp1_2_, 
        temp1_1_, n22}), .B({n20, in3[5:3], n21, in3[1:0]}), .SUM(out2) );
  add_14_DW01_add_3 add_31 ( .A({temp1_6_, n24, temp1_4_, temp1_3_, temp1_2_, 
        temp1_1_, n22}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_14_DW01_add_4 add_30 ( .A({in2[6:4], n23, in2[2], n19, in2[0]}), .B({n20, 
        in3[5:3], n21, in3[1:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_14_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX3 U1 ( .A(in2[1]), .Y(n19) );
  CLKBUFX1TH U2 ( .A(in3[6]), .Y(n20) );
  CLKBUFX40 U3 ( .A(in3[2]), .Y(n21) );
  CLKBUFX40 U4 ( .A(temp1_0_), .Y(n22) );
  CLKBUFX40 U5 ( .A(in2[3]), .Y(n23) );
  CLKBUFX40 U6 ( .A(temp1_5_), .Y(n24) );
endmodule


module tc_sm_59 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  CLKBUFX2TH U3 ( .A(in[6]), .Y(out[4]) );
  NOR3X1TH U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U5 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U6 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U7 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U8 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n28) );
  INVXLTH U12 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n29) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_58 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n23, n24, n25, n26;

  OAI211X1 U3 ( .A0(in[6]), .A1(n24), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI221X2TH U4 ( .A0(n23), .A1(n8), .B0(in[6]), .B1(n25), .C0(n6), .Y(out[2])
         );
  OAI21X1TH U5 ( .A0(n7), .A1(n24), .B0(in[6]), .Y(n5) );
  OAI2B11X4TH U6 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OAI221X1 U7 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n26), .C0(n6), .Y(out[1])
         );
  INVX1 U8 ( .A(in[6]), .Y(n23) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  AOI2BB1X4 U10 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  NAND2BXLTH U11 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  XOR2XLTH U12 ( .A(in[0]), .B(n26), .Y(n10) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U14 ( .A(in[3]), .Y(n24) );
  AOI21X8 U15 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n6) );
  INVXLTH U16 ( .A(in[1]), .Y(n26) );
  INVXLTH U17 ( .A(in[2]), .Y(n25) );
  XOR2XLTH U18 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n9) );
endmodule


module tc_sm_57 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n21, n22, n24, n25, n26, n27, n28,
         n29, n31;

  OAI2BB1X2TH U3 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI221XLTH U4 ( .A0(n24), .A1(n10), .B0(n31), .B1(n28), .C0(n22), .Y(out[2])
         );
  CLKINVX16 U5 ( .A(n21), .Y(n22) );
  CLKINVX1TH U6 ( .A(in[3]), .Y(n27) );
  NOR3X1TH U7 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U8 ( .A(in[5]), .Y(n25) );
  CLKBUFX1TH U9 ( .A(n31), .Y(out[4]) );
  OAI221XLTH U10 ( .A0(n24), .A1(n12), .B0(n31), .B1(n29), .C0(n22), .Y(out[1]) );
  INVXLTH U11 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U13 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U15 ( .A(in[2]), .Y(n28) );
  OAI21XLTH U16 ( .A0(n9), .A1(n27), .B0(n31), .Y(n7) );
  INVX6 U17 ( .A(n8), .Y(n21) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n22), .Y(out[0]) );
  INVXLTH U19 ( .A(n31), .Y(n24) );
  OAI211XLTH U20 ( .A0(n31), .A1(n27), .B0(n7), .C0(n22), .Y(out[3]) );
  OAI33X4 U21 ( .A0(in[4]), .A1(n31), .A2(in[5]), .B0(n13), .B1(n25), .B2(n26), 
        .Y(n8) );
  INVXL U22 ( .A(in[4]), .Y(n26) );
  CLKBUFX40 U23 ( .A(in[6]), .Y(n31) );
endmodule


module tc_sm_56 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n22, n23, n25, n26, n27, n29, n30, n31,
         n32, n33, n34;

  OAI221XL U3 ( .A0(n22), .A1(n12), .B0(in[6]), .B1(n27), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U7 ( .A0(n22), .A1(n10), .B0(in[6]), .B1(n26), .C0(n8), .Y(out[2]) );
  OAI211XLTH U8 ( .A0(in[6]), .A1(n25), .B0(n7), .C0(n8), .Y(out[3]) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U10 ( .A(in[3]), .Y(n25) );
  XNOR2XLTH U11 ( .A(n26), .B(n11), .Y(n10) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U13 ( .A(in[2]), .Y(n26) );
  OAI21XLTH U14 ( .A0(n9), .A1(n25), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U17 ( .A(in[1]), .Y(n27) );
  XNOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVX2 U19 ( .A(in[5]), .Y(n23) );
  INVXLTH U20 ( .A(in[6]), .Y(n22) );
  DLY1X1TH U4 ( .A(in[4]), .Y(n29) );
  AOI33X4 U5 ( .A0(n31), .A1(n32), .A2(n23), .B0(n34), .B1(n33), .B2(in[4]), 
        .Y(n30) );
  CLKINVX40 U6 ( .A(n30), .Y(n8) );
  CLKINVX40 U21 ( .A(n29), .Y(n31) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n32) );
  CLKINVX40 U23 ( .A(n23), .Y(n33) );
  AOI21BX4 U24 ( .A0(n25), .A1(n9), .B0N(in[6]), .Y(n34) );
endmodule


module total_3_test_33 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n63, w5_4_, n4, n5, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n60;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_59 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_58 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_57 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_56 sm_tc_4 ( .out(in1), .in(in) );
  add_14 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_59 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_58 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_57 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_56 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n47), .CK(clk), .RN(n5), .Q(
        h) );
  SDFFRQX1TH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n45), .CK(clk), .RN(n4), 
        .Q(up1[2]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up1[4]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n45), .CK(clk), .RN(n4), 
        .Q(up2[3]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n52), .CK(clk), .RN(n5), 
        .Q(n63) );
  SDFFRQX4TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up2[4]) );
  SDFFRQX2 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n5) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n4) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n53), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRX4 up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n49), .CK(clk), .RN(n4), .Q(n54)
         );
  SDFFRX4 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n53), .CK(clk), .RN(n4), 
        .Q(up1[1]) );
  DLY1X1TH U37 ( .A(n46), .Y(n44) );
  INVXLTH U38 ( .A(n46), .Y(n45) );
  DLY1X1TH U39 ( .A(n50), .Y(n46) );
  INVXLTH U40 ( .A(n46), .Y(n47) );
  INVXLTH U41 ( .A(n50), .Y(n48) );
  DLY1X1TH U42 ( .A(test_se), .Y(n49) );
  INVXLTH U43 ( .A(test_se), .Y(n50) );
  INVXLTH U44 ( .A(n44), .Y(n51) );
  INVXLTH U45 ( .A(n44), .Y(n52) );
  INVXLTH U46 ( .A(n46), .Y(n53) );
  CLKINVX40 U47 ( .A(n54), .Y(n60) );
  CLKINVX40 U48 ( .A(n60), .Y(up1[0]) );
  DLY1X1TH U49 ( .A(n63), .Y(up3[3]) );
endmodule


module sm_tc_55 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n17, n18, n21, n22, n23, n24, n25;

  AOI31X1 U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n17), .Y(out[4]) );
  OAI2BB2X1TH U5 ( .B0(n17), .B1(n4), .A0N(in[3]), .A1N(n17), .Y(out[3]) );
  INVX4 U6 ( .A(in[4]), .Y(n17) );
  XNOR2X1 U7 ( .A(n22), .B(n8), .Y(n5) );
  NOR2X4 U8 ( .A(in[1]), .B(n25), .Y(n8) );
  AO21XL U9 ( .A0(n25), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2X4 U10 ( .B0(n17), .B1(n6), .A0N(in[1]), .A1N(n17), .Y(out[1]) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX1TH U12 ( .A(n25), .Y(out[0]) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U14 ( .AN(n6), .B(n25), .Y(n3) );
  INVX2 U16 ( .A(in[2]), .Y(n18) );
  CLKINVX40 U2 ( .A(n18), .Y(n21) );
  CLKINVX40 U4 ( .A(n21), .Y(n22) );
  OAI2BB2X2 U15 ( .B0(n17), .B1(n5), .A0N(n17), .A1N(n23), .Y(out[2]) );
  CLKINVX40 U17 ( .A(n22), .Y(n23) );
  XOR2X1 U18 ( .A(n24), .B(in[3]), .Y(n4) );
  CLKAND2X12 U19 ( .A(n8), .B(n22), .Y(n24) );
  CLKBUFX40 U20 ( .A(in[0]), .Y(n25) );
endmodule


module sm_tc_54 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n17, n18, n22, n23, n25, n26;

  CLKBUFX1 U3 ( .A(out[4]), .Y(out[5]) );
  BUFX2 U4 ( .A(in[4]), .Y(n18) );
  NOR2X2TH U5 ( .A(in[1]), .B(n17), .Y(n8) );
  INVX4 U6 ( .A(n18), .Y(n22) );
  BUFX10 U7 ( .A(in[0]), .Y(n17) );
  OAI2BB2X1TH U8 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U9 ( .A(n17), .Y(out[0]) );
  AO21X2TH U10 ( .A0(n17), .A1(in[1]), .B0(n8), .Y(n6) );
  AOI31X2TH U11 ( .A0(n3), .A1(n4), .A2(n25), .B0(n22), .Y(out[4]) );
  OAI2BB2X2 U12 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  OAI22X2 U13 ( .A0(n18), .A1(n23), .B0(n22), .B1(n25), .Y(out[2]) );
  INVX2TH U14 ( .A(in[2]), .Y(n23) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[6]) );
  NOR2BXLTH U17 ( .AN(n6), .B(n17), .Y(n3) );
  XNOR2X1TH U18 ( .A(n23), .B(n8), .Y(n5) );
  CLKBUFX40 U2 ( .A(n5), .Y(n25) );
  XOR2X1 U16 ( .A(n26), .B(in[3]), .Y(n4) );
  CLKAND2X12 U19 ( .A(n8), .B(n23), .Y(n26) );
endmodule


module sm_tc_53 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n27, n28, n30, n33, n34;

  NOR2X4 U2 ( .A(n28), .B(in[0]), .Y(n8) );
  BUFX6 U3 ( .A(in[4]), .Y(n27) );
  XNOR2X1 U4 ( .A(n34), .B(n8), .Y(n5) );
  INVX4TH U5 ( .A(n27), .Y(n33) );
  OAI2BB2X1TH U6 ( .B0(n33), .B1(n6), .A0N(n28), .A1N(n33), .Y(out[1]) );
  CLKBUFX2TH U7 ( .A(in[1]), .Y(n28) );
  AOI31X2TH U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n33), .Y(out[4]) );
  AO21X2 U9 ( .A0(in[0]), .A1(n28), .B0(n8), .Y(n6) );
  CLKBUFX2 U10 ( .A(in[0]), .Y(out[0]) );
  OAI22X2 U11 ( .A0(n27), .A1(n34), .B0(n33), .B1(n5), .Y(out[2]) );
  OAI2BB2X4TH U12 ( .B0(n33), .B1(n4), .A0N(in[3]), .A1N(n33), .Y(out[3]) );
  INVXLTH U13 ( .A(n30), .Y(out[5]) );
  INVX2TH U14 ( .A(in[2]), .Y(n34) );
  XNOR2X2TH U15 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKNAND2X2 U16 ( .A(n8), .B(n34), .Y(n7) );
  INVXLTH U17 ( .A(n30), .Y(out[6]) );
  NOR2BXLTH U18 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U19 ( .A(out[4]), .Y(n30) );
endmodule


module sm_tc_52 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n18, n19, n20, n24, n25;

  CLKBUFX1TH U2 ( .A(out[6]), .Y(out[5]) );
  AOI31X4 U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n25), .Y(out[6]) );
  XNOR2X1 U4 ( .A(n24), .B(n8), .Y(n5) );
  NAND2X6 U5 ( .A(n19), .B(n20), .Y(n4) );
  CLKNAND2X2 U6 ( .A(n7), .B(in[3]), .Y(n19) );
  INVXLTH U7 ( .A(n7), .Y(n17) );
  OAI2BB2X1TH U8 ( .B0(n25), .B1(n4), .A0N(in[3]), .A1N(n25), .Y(out[3]) );
  OAI22X1TH U9 ( .A0(in[4]), .A1(n24), .B0(n25), .B1(n5), .Y(out[2]) );
  CLKBUFX1TH U10 ( .A(in[0]), .Y(out[0]) );
  NOR2X2TH U11 ( .A(in[1]), .B(in[0]), .Y(n8) );
  NAND2X4 U12 ( .A(n17), .B(n18), .Y(n20) );
  INVXLTH U13 ( .A(in[3]), .Y(n18) );
  NOR2BX1TH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX1TH U15 ( .A(in[2]), .Y(n24) );
  CLKINVX2TH U16 ( .A(in[4]), .Y(n25) );
  NAND2XLTH U17 ( .A(n8), .B(n24), .Y(n7) );
  CLKBUFX1TH U18 ( .A(out[6]), .Y(out[4]) );
  OAI2BB2X2 U19 ( .B0(n25), .B1(n6), .A0N(in[1]), .A1N(n25), .Y(out[1]) );
  AO21XLTH U20 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_13_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X4TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_13_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, n1;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry_6_), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry_2_), .S(SUM[1]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_13_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, n1, n2;

  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry_2_), .S(SUM[1]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry_6_), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_13_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_13_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   carry_4_, carry_3_, carry_2_, n1, n2, n3, n4, n5, n6;
  wire   [6:5] carry;

  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX4 U1_2 ( .A(B[2]), .B(carry_2_), .CI(A[2]), .CO(carry_3_), .S(SUM[2])
         );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHX2 U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry_2_), .S(SUM[1]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry[5]), .S(SUM[4])
         );
  XOR2X2 U1 ( .A(n2), .B(carry_3_), .Y(SUM[3]) );
  NAND2XLTH U4 ( .A(A[3]), .B(B[3]), .Y(n5) );
  NAND2XLTH U5 ( .A(carry_3_), .B(B[3]), .Y(n4) );
  NAND3X2 U6 ( .A(n3), .B(n4), .C(n5), .Y(carry_4_) );
  NAND2XLTH U7 ( .A(carry_3_), .B(A[3]), .Y(n3) );
  AND2XLTH U8 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR2X1 U3 ( .A(n6), .B(A[3]), .Y(n2) );
  CLKINVX40 U9 ( .A(B[3]), .Y(n6) );
endmodule


module add_13_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n3, n1;
  wire   [6:2] carry;

  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(n3) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKBUFX40 U3 ( .A(n3), .Y(SUM[2]) );
endmodule


module add_13 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;

  add_13_DW01_add_0 add_34 ( .A({temp1_6_, n28, n27, temp1_3_, temp1_2_, 
        temp1_1_, n30}), .B({in2[6:4], n23, n29, n21, in2[0]}), .SUM(out3) );
  add_13_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, n20, temp2_2_, 
        temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_13_DW01_add_2 add_32 ( .A({temp1_6_, n28, n27, temp1_3_, temp1_2_, 
        temp1_1_, n30}), .B({in3[6:3], n26, in3[1], n24}), .SUM(out2) );
  add_13_DW01_add_3 add_31 ( .A({temp1_6_, n28, n27, temp1_3_, temp1_2_, 
        temp1_1_, n30}), .B({temp2_6_, temp2_5_, temp2_4_, n20, temp2_2_, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_13_DW01_add_4 add_30 ( .A({in2[6:4], n23, n29, n21, in2[0]}), .B({
        in3[6:3], n26, in3[1], n24}), .SUM({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_13_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  INVX4 U1 ( .A(n22), .Y(n23) );
  CLKINVX12 U2 ( .A(temp2_3_), .Y(n19) );
  INVX12 U3 ( .A(n19), .Y(n20) );
  BUFX3 U4 ( .A(in2[1]), .Y(n21) );
  CLKBUFX1TH U5 ( .A(in3[0]), .Y(n24) );
  CLKINVX1TH U6 ( .A(n25), .Y(n26) );
  INVX2TH U13 ( .A(in3[2]), .Y(n25) );
  CLKINVX6 U14 ( .A(in2[3]), .Y(n22) );
  CLKBUFX40 U15 ( .A(temp1_4_), .Y(n27) );
  CLKBUFX40 U16 ( .A(temp1_5_), .Y(n28) );
  CLKBUFX40 U17 ( .A(in2[2]), .Y(n29) );
  CLKBUFX40 U18 ( .A(temp1_0_), .Y(n30) );
endmodule


module tc_sm_55 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U10 ( .A(in[4]), .Y(n28) );
  INVXLTH U11 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI2BB1XLTH U19 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI211XLTH U20 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
endmodule


module tc_sm_54 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n6, n14, n16, n17, n18, n19, n20;

  OAI2BB1X2 U3 ( .A0N(n18), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI2B11X2 U4 ( .A1N(n14), .A0(n18), .B0(n7), .C0(n6), .Y(out[3]) );
  INVX1 U5 ( .A(in[6]), .Y(n14) );
  OAI221X1 U6 ( .A0(n14), .A1(n10), .B0(in[6]), .B1(n19), .C0(n6), .Y(out[2])
         );
  CLKINVX1TH U7 ( .A(in[3]), .Y(n18) );
  BUFX10 U8 ( .A(n8), .Y(n6) );
  NAND2BXLTH U9 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  OAI221XLTH U10 ( .A0(n14), .A1(n12), .B0(in[6]), .B1(n20), .C0(n6), .Y(
        out[1]) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U13 ( .A(in[1]), .Y(n20) );
  XNOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U15 ( .A(n19), .B(n11), .Y(n10) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U17 ( .A(in[2]), .Y(n19) );
  OAI21XLTH U18 ( .A0(n9), .A1(n18), .B0(in[6]), .Y(n7) );
  INVX2 U19 ( .A(in[5]), .Y(n16) );
  OAI33X4 U20 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n16), .B2(
        n17), .Y(n8) );
  INVXL U21 ( .A(in[4]), .Y(n17) );
endmodule


module tc_sm_53 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n21,
         n22;

  OAI221XL U3 ( .A0(n14), .A1(n10), .B0(in[6]), .B1(n18), .C0(n22), .Y(out[2])
         );
  OAI221XL U4 ( .A0(n14), .A1(n12), .B0(in[6]), .B1(n19), .C0(n22), .Y(out[1])
         );
  OAI211XL U5 ( .A0(in[6]), .A1(n17), .B0(n7), .C0(n22), .Y(out[3]) );
  OAI2BB1X4 U6 ( .A0N(n17), .A1N(n9), .B0(in[6]), .Y(n13) );
  INVXLTH U7 ( .A(in[6]), .Y(n14) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n17) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U10 ( .A(in[1]), .Y(n19) );
  XNOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U12 ( .A(n18), .B(n11), .Y(n10) );
  NOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U14 ( .A(in[2]), .Y(n18) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U16 ( .A0(n9), .A1(n17), .B0(in[6]), .Y(n7) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n22), .Y(out[0]) );
  OAI33X4 U18 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n15), .B2(
        n16), .Y(n8) );
  INVXL U19 ( .A(in[5]), .Y(n15) );
  INVXL U20 ( .A(in[4]), .Y(n16) );
  CLKINVX40 U21 ( .A(n8), .Y(n21) );
  CLKINVX40 U22 ( .A(n21), .Y(n22) );
endmodule


module tc_sm_52 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n22, n23, n24, n25;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  AOI21X6 U3 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n6) );
  AOI2BB1X2 U4 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  OAI221XL U5 ( .A0(n22), .A1(n8), .B0(in[6]), .B1(n24), .C0(n6), .Y(out[2])
         );
  INVXLTH U6 ( .A(in[6]), .Y(n22) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U9 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U10 ( .A(in[2]), .Y(n24) );
  XOR2XLTH U11 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n9) );
  XOR2XLTH U13 ( .A(in[0]), .B(n25), .Y(n10) );
  INVXLTH U14 ( .A(in[1]), .Y(n25) );
  OAI21XLTH U15 ( .A0(n7), .A1(n23), .B0(in[6]), .Y(n5) );
  INVXLTH U16 ( .A(in[3]), .Y(n23) );
  OAI221XLTH U17 ( .A0(n22), .A1(n10), .B0(in[6]), .B1(n25), .C0(n6), .Y(
        out[1]) );
  OAI211XLTH U18 ( .A0(in[6]), .A1(n23), .B0(n5), .C0(n6), .Y(out[3]) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n6), .Y(out[0]) );
endmodule


module total_3_test_34 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n53, w5_4_, n4, n5, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_55 sm_tc_1 ( .out(a1), .in({a[4], n40, a[2:0]}) );
  sm_tc_54 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_53 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_52 sm_tc_4 ( .out(in1), .in(in) );
  add_13 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_55 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_54 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_53 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_52 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n46), .CK(clk), .RN(n4), 
        .Q(up3[3]) );
  SDFFRQXLTH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n45), .CK(clk), .RN(n5), .Q(
        h) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n49), .CK(clk), .RN(n4), .Q(
        up1[0]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n41), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n46), .CK(clk), .RN(n4), 
        .Q(up2[3]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n41), .CK(clk), .RN(n5), 
        .Q(up1[2]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n42), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n42), .CK(clk), .RN(n4), 
        .Q(n53) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRQX2 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n45), .CK(clk), .RN(n4), 
        .Q(up1[1]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n5) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n4) );
  CLKBUFX40 U37 ( .A(a[3]), .Y(n40) );
  INVXLTH U38 ( .A(n44), .Y(n41) );
  INVXLTH U39 ( .A(n43), .Y(n42) );
  DLY1X1TH U40 ( .A(n47), .Y(n43) );
  DLY1X1TH U41 ( .A(n47), .Y(n44) );
  INVXLTH U42 ( .A(n44), .Y(n45) );
  INVXLTH U43 ( .A(n43), .Y(n46) );
  INVXLTH U44 ( .A(test_se), .Y(n47) );
  INVXLTH U45 ( .A(n44), .Y(n48) );
  INVXLTH U46 ( .A(n43), .Y(n49) );
  INVXLTH U47 ( .A(n44), .Y(n50) );
  INVXLTH U48 ( .A(n43), .Y(n51) );
  DLY1X1TH U49 ( .A(n53), .Y(up2[2]) );
endmodule


module sm_tc_51 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n23;

  AOI31X1 U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  OAI22XLTH U3 ( .A0(in[4]), .A1(n23), .B0(n22), .B1(n5), .Y(out[2]) );
  XNOR2X1 U4 ( .A(n23), .B(n8), .Y(n5) );
  CLKBUFX4 U5 ( .A(in[0]), .Y(out[0]) );
  NOR2X6 U6 ( .A(in[1]), .B(out[0]), .Y(n8) );
  AO21X1 U7 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  INVX3TH U8 ( .A(in[4]), .Y(n22) );
  XNOR2X1TH U9 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X2 U10 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  OAI2BB2X1TH U11 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  INVX1TH U12 ( .A(in[2]), .Y(n23) );
  NAND2XLTH U13 ( .A(n8), .B(n23), .Y(n7) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U16 ( .AN(n6), .B(out[0]), .Y(n3) );
endmodule


module sm_tc_50 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n27, n3, n4, n5, n6, n7, n8, n17, n21, n22, n26;

  AOI31X2 U2 ( .A0(n3), .A1(n5), .A2(n4), .B0(n21), .Y(n27) );
  BUFX4 U3 ( .A(in[4]), .Y(n17) );
  BUFX2TH U4 ( .A(out[4]), .Y(out[5]) );
  XNOR2X1TH U5 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U6 ( .A(n8), .B(n26), .Y(n7) );
  XNOR2X1 U7 ( .A(n26), .B(n8), .Y(n5) );
  OAI2BB2X1 U8 ( .B0(n21), .B1(n4), .A0N(in[3]), .A1N(n21), .Y(out[3]) );
  OAI22XLTH U9 ( .A0(n17), .A1(n26), .B0(n21), .B1(n5), .Y(out[2]) );
  OAI2BB2X2 U10 ( .B0(n21), .B1(n6), .A0N(in[1]), .A1N(n21), .Y(out[1]) );
  INVX3TH U11 ( .A(n17), .Y(n21) );
  NOR2X3 U12 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[6]) );
  AO21XLTH U14 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKINVX1TH U15 ( .A(in[2]), .Y(n22) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  BUFX2TH U17 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX40 U18 ( .A(n27), .Y(out[4]) );
  CLKBUFX40 U19 ( .A(n22), .Y(n26) );
endmodule


module sm_tc_49 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n35, n36, n39, n40, n41, n42;

  OAI2BB2X4 U2 ( .B0(n40), .B1(n6), .A0N(n40), .A1N(in[1]), .Y(out[1]) );
  NOR2X2 U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X1TH U4 ( .A(n36), .B(n41), .Y(n5) );
  XNOR2X1TH U5 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U6 ( .A(n41), .B(n36), .Y(n7) );
  AO21XLTH U7 ( .A0(in[0]), .A1(in[1]), .B0(n41), .Y(n6) );
  CLKBUFX1TH U8 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U9 ( .A(out[5]), .Y(out[6]) );
  BUFX2TH U10 ( .A(out[5]), .Y(out[4]) );
  AOI31X4 U11 ( .A0(n3), .A1(n4), .A2(n42), .B0(n40), .Y(out[5]) );
  CLKINVX1TH U12 ( .A(in[2]), .Y(n36) );
  INVX4TH U13 ( .A(in[4]), .Y(n35) );
  OAI22X4TH U14 ( .A0(in[4]), .A1(n36), .B0(n40), .B1(n42), .Y(out[2]) );
  OAI2BB2X1TH U15 ( .B0(n40), .B1(n4), .A0N(in[3]), .A1N(n40), .Y(out[3]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKINVX40 U17 ( .A(n35), .Y(n39) );
  CLKINVX40 U18 ( .A(n39), .Y(n40) );
  CLKBUFX40 U19 ( .A(n8), .Y(n41) );
  CLKBUFX40 U20 ( .A(n5), .Y(n42) );
endmodule


module sm_tc_48 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  XNOR2X1 U2 ( .A(n7), .B(in[3]), .Y(n4) );
  NOR2X2TH U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVXLTH U4 ( .A(out[4]), .Y(n18) );
  OAI2BB2X1TH U5 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  AOI31X2TH U6 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  CLKINVX1TH U7 ( .A(in[2]), .Y(n21) );
  CLKINVX2TH U8 ( .A(in[4]), .Y(n22) );
  NOR2BXLTH U9 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U10 ( .A(n18), .Y(out[5]) );
  OAI22X1TH U11 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  OAI2BB2X1TH U12 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U13 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U14 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U15 ( .A(n21), .B(n8), .Y(n5) );
  NAND2XLTH U16 ( .A(n8), .B(n21), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_12_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X4 U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  XOR2X2TH U2 ( .A(B[6]), .B(A[6]), .Y(n2) );
  AND2XLTH U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_12_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR2X1 U3 ( .A(A[6]), .B(n3), .Y(n2) );
  CLKXOR2X8 U4 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  CLKINVX40 U5 ( .A(B[6]), .Y(n3) );
endmodule


module add_12_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_12_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR3X2 U3 ( .A(A[6]), .B(n3), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
  CLKINVX40 U5 ( .A(B[6]), .Y(n3) );
endmodule


module add_12_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;
  wire   [6:2] carry;

  NAND3X2 U11 ( .A(n2), .B(n3), .C(n4), .Y(carry[6]) );
  NAND2X2 U13 ( .A(A[2]), .B(B[2]), .Y(n9) );
  ADDFHX2 U1_3 ( .A(A[3]), .B(carry[3]), .CI(B[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_1 ( .A(n5), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND2X4 U1 ( .A(n12), .B(n13), .Y(SUM[5]) );
  INVX2TH U2 ( .A(n1), .Y(n10) );
  XNOR2X2 U3 ( .A(n14), .B(carry[2]), .Y(SUM[2]) );
  NAND2X2 U4 ( .A(carry[2]), .B(B[2]), .Y(n8) );
  CLKNAND2X4 U7 ( .A(n10), .B(carry[5]), .Y(n13) );
  XOR2X1TH U8 ( .A(A[5]), .B(B[5]), .Y(n1) );
  NAND2X2 U9 ( .A(n1), .B(n11), .Y(n12) );
  INVXLTH U10 ( .A(carry[5]), .Y(n11) );
  CLKNAND2X2 U12 ( .A(B[5]), .B(A[5]), .Y(n4) );
  XNOR2X4TH U14 ( .A(B[2]), .B(A[2]), .Y(n14) );
  CLKNAND2X2 U15 ( .A(carry[5]), .B(A[5]), .Y(n3) );
  AND2XLTH U16 ( .A(B[0]), .B(A[0]), .Y(n5) );
  CLKXOR2X1TH U17 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND3X4 U18 ( .A(n7), .B(n8), .C(n9), .Y(carry[3]) );
  AND2X8 U5 ( .A(carry[2]), .B(A[2]), .Y(n15) );
  CLKINVX40 U6 ( .A(n15), .Y(n7) );
  AND2X8 U19 ( .A(carry[5]), .B(B[5]), .Y(n16) );
  CLKINVX40 U20 ( .A(n16), .Y(n2) );
endmodule


module add_12_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X2 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_12 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n18, n19, n20, n21, n22, n23, n24, n25, n26;

  add_12_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in2[6:5], n20, in2[3], n26, 
        in2[1:0]}), .SUM(out3) );
  add_12_DW01_add_1 add_33 ( .A({temp2_6_, n19, temp2_4_, temp2_3_, n18, 
        temp2_1_, temp2_0_}), .B({n24, in[5:0]}), .SUM(out1) );
  add_12_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in3[6:3], n25, in3[1], n22}), 
        .SUM(out2) );
  add_12_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({temp2_6_, n19, temp2_4_, temp2_3_, 
        n18, temp2_1_, temp2_0_}), .SUM(out) );
  add_12_DW01_add_4 add_30 ( .A({in2[6:5], n20, in2[3], n26, in2[1:0]}), .B({
        in3[6:3], n25, in3[1], n22}), .SUM({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_12_DW01_add_5 add_29 ( .A({n23, in[5:0]}), .B(in1), .SUM({temp1_6_, 
        temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2TH U1 ( .A(temp2_5_), .Y(n19) );
  BUFX2 U2 ( .A(in2[2]), .Y(n21) );
  BUFX8 U3 ( .A(temp2_2_), .Y(n18) );
  CLKBUFX1TH U4 ( .A(in2[4]), .Y(n20) );
  CLKBUFX40 U5 ( .A(in3[0]), .Y(n22) );
  DLY1X1TH U6 ( .A(in[6]), .Y(n23) );
  DLY1X1TH U13 ( .A(in[6]), .Y(n24) );
  CLKBUFX40 U14 ( .A(in3[2]), .Y(n25) );
  CLKBUFX40 U15 ( .A(n21), .Y(n26) );
endmodule


module tc_sm_51 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(in[6]), .Y(n26) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n28) );
  INVXLTH U12 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_50 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n20, n21, n22, n23, n24, n25, n28,
         n29, n30, n31, n32, n33, n35, n36, n37, n38, n39;

  OAI2BB1X4 U3 ( .A0N(n31), .A1N(n9), .B0(in[6]), .Y(n13) );
  OA21XL U4 ( .A0(n36), .A1(n31), .B0(n7), .Y(n20) );
  NAND2XLTH U5 ( .A(n20), .B(n21), .Y(out[3]) );
  NAND3XL U6 ( .A(n22), .B(n23), .C(n21), .Y(out[1]) );
  OR2X2 U7 ( .A(n39), .B(n12), .Y(n22) );
  OR3X1 U8 ( .A(n24), .B(n25), .C(n38), .Y(out[2]) );
  NOR2XL U9 ( .A(n28), .B(n10), .Y(n24) );
  BUFX10 U10 ( .A(n8), .Y(n21) );
  NAND2BX2TH U12 ( .AN(in[0]), .B(n35), .Y(out[0]) );
  OR2XLTH U13 ( .A(n36), .B(n33), .Y(n23) );
  NOR2XLTH U14 ( .A(n36), .B(n32), .Y(n25) );
  XNOR2X1TH U15 ( .A(n32), .B(n11), .Y(n10) );
  OAI33X4 U16 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n29), .B2(
        n30), .Y(n8) );
  INVXLTH U17 ( .A(n36), .Y(n28) );
  CLKINVX1TH U18 ( .A(in[3]), .Y(n31) );
  NOR3X1TH U19 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U20 ( .A(in[4]), .Y(n30) );
  INVXLTH U21 ( .A(in[5]), .Y(n29) );
  INVXLTH U22 ( .A(in[1]), .Y(n33) );
  XNOR2XLTH U23 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U24 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U25 ( .A(in[2]), .Y(n32) );
  CLKBUFX1TH U27 ( .A(n36), .Y(out[4]) );
  CLKINVX40 U11 ( .A(n38), .Y(n35) );
  CLKBUFX40 U26 ( .A(in[6]), .Y(n36) );
  OA21X4 U28 ( .A0(n9), .A1(n31), .B0(in[6]), .Y(n37) );
  CLKINVX40 U29 ( .A(n37), .Y(n7) );
  CLKINVX40 U30 ( .A(n21), .Y(n38) );
  INVXLTH U31 ( .A(in[6]), .Y(n39) );
endmodule


module tc_sm_49 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n26, n27,
         n28;

  NAND2BX2 U3 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211X2 U4 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221X2 U5 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1])
         );
  OAI221X2 U6 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2])
         );
  INVXLTH U7 ( .A(in[6]), .Y(n19) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n22) );
  XNOR2XLTH U10 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U12 ( .A(in[2]), .Y(n23) );
  OAI21XLTH U13 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  INVXLTH U14 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n12) );
  CLKBUFX1TH U16 ( .A(in[6]), .Y(out[4]) );
  INVX2 U18 ( .A(in[5]), .Y(n20) );
  INVXL U20 ( .A(in[4]), .Y(n21) );
  AOI33X4 U17 ( .A0(n21), .A1(n27), .A2(n20), .B0(n28), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U19 ( .A(n26), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n27) );
  AOI21BX4 U22 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n28) );
endmodule


module tc_sm_48 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n26, n27, n28,
         n29;

  OAI221XL U3 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n29), .Y(out[2])
         );
  OAI221XL U4 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n29), .Y(out[1])
         );
  OAI211XL U5 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n29), .Y(out[3]) );
  INVXLTH U6 ( .A(in[4]), .Y(n21) );
  CLKINVX1TH U7 ( .A(in[3]), .Y(n22) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  NAND2BXLTH U10 ( .AN(in[0]), .B(n29), .Y(out[0]) );
  INVXLTH U11 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U13 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U16 ( .A(in[2]), .Y(n23) );
  OAI21XLTH U17 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  INVXLTH U18 ( .A(in[6]), .Y(n19) );
  INVX2 U19 ( .A(in[5]), .Y(n20) );
  AOI33X4 U8 ( .A0(n21), .A1(n27), .A2(n20), .B0(n28), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U20 ( .A(in[6]), .Y(n27) );
  AOI21BX4 U21 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n28) );
  CLKINVX40 U22 ( .A(n26), .Y(n29) );
endmodule


module total_3_test_35 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n66, n67, w5_4_, n4, n5, n6, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_51 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_50 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_49 sm_tc_3 ( .out(c1), .in({n4, c[3:0]}) );
  sm_tc_48 sm_tc_4 ( .out(in1), .in(in) );
  add_12 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3({c1[6:4], n46, c1[2:0]}), .in(in1) );
  tc_sm_51 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_50 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_49 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_48 tc_sm_4 ( .out(w8), .in({n58, w88[5:0]}) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n57), .CK(clk), .RN(n5), 
        .Q(up3[3]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n47), .CK(clk), .RN(n5), 
        .Q(n67) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n52), .CK(clk), .RN(n6), .Q(
        h) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n56), .CK(clk), .RN(n5), .Q(
        up1[0]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n57), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n47), .CK(clk), .RN(n5), 
        .Q(n66) );
  SDFFRQXLTH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n56), .CK(clk), .RN(n5), 
        .Q(up2[1]) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n54), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQX1TH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n54), .CK(clk), .RN(n5), 
        .Q(up2[2]) );
  CLKBUFX1TH U3 ( .A(c[4]), .Y(n4) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n5) );
  CLKBUFX1TH U5 ( .A(rst), .Y(n6) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n55), .CK(clk), .RN(n5), 
        .Q(up1[3]) );
  SDFFRX4 up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n55), .CK(clk), .RN(n6), 
        .Q(up1[4]) );
  SDFFRHQX8 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n52), .CK(clk), .RN(n6), 
        .Q(up1[2]) );
  SDFFRX4 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  CLKBUFX40 U38 ( .A(c1[3]), .Y(n46) );
  INVXLTH U39 ( .A(n50), .Y(n47) );
  INVXLTH U40 ( .A(n49), .Y(n48) );
  DLY1X1TH U41 ( .A(n53), .Y(n49) );
  DLY1X1TH U42 ( .A(n53), .Y(n50) );
  INVXLTH U43 ( .A(n50), .Y(n51) );
  INVXLTH U44 ( .A(n49), .Y(n52) );
  INVXLTH U45 ( .A(test_se), .Y(n53) );
  INVXLTH U46 ( .A(n50), .Y(n54) );
  INVXLTH U47 ( .A(n49), .Y(n55) );
  INVXLTH U48 ( .A(n50), .Y(n56) );
  INVXLTH U49 ( .A(n49), .Y(n57) );
  CLKBUFX40 U50 ( .A(w88[6]), .Y(n58) );
  DLY1X1TH U51 ( .A(n66), .Y(up2[3]) );
  DLY1X1TH U52 ( .A(n67), .Y(up3[4]) );
endmodule


module sm_tc_47 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n17, n18, n22, n23, n26;

  AO21X1 U2 ( .A0(n18), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X8 U3 ( .A(in[1]), .B(n18), .Y(n8) );
  BUFX10 U4 ( .A(in[4]), .Y(n17) );
  INVX5TH U5 ( .A(n17), .Y(n22) );
  BUFX10 U6 ( .A(in[0]), .Y(n18) );
  XNOR2X2TH U7 ( .A(n23), .B(n8), .Y(n5) );
  BUFX2TH U8 ( .A(n18), .Y(out[0]) );
  INVX2 U10 ( .A(in[2]), .Y(n23) );
  OAI2BB2XLTH U11 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X4 U13 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  AOI31X2TH U15 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U16 ( .AN(n6), .B(n18), .Y(n3) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[5]) );
  OAI22XLTH U18 ( .A0(n17), .A1(n23), .B0(n22), .B1(n5), .Y(out[2]) );
  XOR2X1 U9 ( .A(n26), .B(in[3]), .Y(n4) );
  CLKAND2X12 U14 ( .A(n8), .B(n23), .Y(n26) );
endmodule


module sm_tc_46 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n24, n25, n28, n29, n30;

  OAI22X1 U2 ( .A0(in[4]), .A1(n25), .B0(n24), .B1(n5), .Y(out[2]) );
  INVX2 U5 ( .A(in[2]), .Y(n25) );
  OAI2BB2X1 U6 ( .B0(n24), .B1(n4), .A0N(in[3]), .A1N(n24), .Y(out[3]) );
  INVX2TH U7 ( .A(in[4]), .Y(n24) );
  CLKBUFX2TH U9 ( .A(in[0]), .Y(out[0]) );
  AO21X2 U10 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X2 U12 ( .B0(n24), .B1(n6), .A0N(in[1]), .A1N(n24), .Y(out[1]) );
  AOI31X2TH U14 ( .A0(n3), .A1(n4), .A2(n5), .B0(n24), .Y(out[4]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  XOR2X1 U3 ( .A(n25), .B(n28), .Y(n5) );
  CLKINVX40 U4 ( .A(n8), .Y(n28) );
  OR2X8 U8 ( .A(in[1]), .B(in[0]), .Y(n29) );
  CLKINVX40 U13 ( .A(n29), .Y(n8) );
  XOR2X1 U17 ( .A(n30), .B(in[3]), .Y(n4) );
  CLKAND2X12 U18 ( .A(n8), .B(n25), .Y(n30) );
endmodule


module sm_tc_45 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n24, n25, n26, n30, n31, n34;

  CLKBUFX4 U2 ( .A(in[1]), .Y(n26) );
  OAI22X4 U4 ( .A0(n25), .A1(n31), .B0(n30), .B1(n5), .Y(out[2]) );
  NOR2X4 U7 ( .A(n26), .B(in[0]), .Y(n8) );
  BUFX2TH U8 ( .A(in[4]), .Y(n25) );
  INVX2 U9 ( .A(n25), .Y(n30) );
  XNOR2X1 U10 ( .A(n31), .B(n8), .Y(n5) );
  INVX2 U11 ( .A(in[2]), .Y(n31) );
  AND2X1TH U12 ( .A(in[0]), .B(n26), .Y(n24) );
  OR2X1 U13 ( .A(n24), .B(n8), .Y(n6) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX1TH U16 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[5]) );
  AOI31X2TH U18 ( .A0(n3), .A1(n4), .A2(n5), .B0(n30), .Y(out[4]) );
  NOR2BXLTH U19 ( .AN(n6), .B(in[0]), .Y(n3) );
  AO2B2X4 U3 ( .B0(in[3]), .B1(n30), .A0(n25), .A1N(n4), .Y(out[3]) );
  AO2B2BX4 U5 ( .A0(n25), .A1N(n6), .B0(n26), .B1N(n25), .Y(out[1]) );
  XOR2X1 U6 ( .A(n34), .B(in[3]), .Y(n4) );
  CLKAND2X12 U14 ( .A(n8), .B(n31), .Y(n34) );
endmodule


module sm_tc_44 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  AOI31X4 U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  XNOR2X2TH U3 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI22X1TH U4 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  BUFX2 U5 ( .A(in[0]), .Y(out[0]) );
  XNOR2X1 U6 ( .A(n21), .B(n8), .Y(n5) );
  NOR2X2TH U7 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U8 ( .A(in[2]), .Y(n21) );
  OAI2BB2X4TH U9 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKINVX2TH U10 ( .A(in[4]), .Y(n22) );
  INVXLTH U11 ( .A(out[4]), .Y(n18) );
  INVXLTH U12 ( .A(n18), .Y(out[5]) );
  INVXLTH U13 ( .A(n18), .Y(out[6]) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2BB2X1TH U15 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  NAND2XLTH U16 ( .A(n8), .B(n21), .Y(n7) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_11_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_11_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [6:2] carry;

  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR2XL U1 ( .A(B[4]), .B(A[4]), .Y(n5) );
  CLKNAND2X4 U2 ( .A(A[4]), .B(B[4]), .Y(n8) );
  NAND2X1 U3 ( .A(n9), .B(B[4]), .Y(n7) );
  AND2X1TH U5 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X2 U6 ( .A(n5), .B(n9), .Y(SUM[4]) );
  NAND3X2TH U7 ( .A(n6), .B(n7), .C(n8), .Y(carry[5]) );
  XOR3X1TH U8 ( .A(A[1]), .B(n1), .C(B[1]), .Y(SUM[1]) );
  CLKXOR2X1TH U9 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND3X2TH U10 ( .A(n3), .B(n2), .C(n4), .Y(carry[2]) );
  NAND2XLTH U11 ( .A(n1), .B(B[1]), .Y(n4) );
  NAND2XLTH U12 ( .A(A[1]), .B(n1), .Y(n2) );
  NAND2XLTH U13 ( .A(A[1]), .B(B[1]), .Y(n3) );
  CLKBUFX40 U4 ( .A(carry[4]), .Y(n9) );
  AND2X8 U14 ( .A(n9), .B(A[4]), .Y(n10) );
  CLKINVX40 U15 ( .A(n10), .Y(n6) );
endmodule


module add_11_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_11_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3XL U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_11_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X3 U1 ( .A(A[2]), .B(B[2]), .Y(n2) );
  XOR2X1 U2 ( .A(n2), .B(carry[2]), .Y(SUM[2]) );
  NAND2X1 U3 ( .A(carry[2]), .B(B[2]), .Y(n3) );
  NAND2X1 U4 ( .A(carry[2]), .B(A[2]), .Y(n4) );
  NAND2X1 U5 ( .A(B[2]), .B(A[2]), .Y(n5) );
  NAND3X4 U6 ( .A(n3), .B(n4), .C(n5), .Y(carry[3]) );
  CLKXOR2X2TH U7 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U8 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_11_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [6:2] carry;

  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(carry[3]), .CI(B[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  NAND2XLTH U2 ( .A(n7), .B(n3), .Y(n4) );
  INVXL U4 ( .A(n7), .Y(n2) );
  INVXLTH U5 ( .A(A[0]), .Y(n3) );
  AND2XLTH U6 ( .A(n7), .B(A[0]), .Y(n1) );
  AND2X8 U1 ( .A(n4), .B(n5), .Y(n6) );
  CLKINVX40 U3 ( .A(n6), .Y(SUM[0]) );
  CLKBUFX40 U7 ( .A(B[0]), .Y(n7) );
  AND2X8 U8 ( .A(n2), .B(A[0]), .Y(n8) );
  CLKINVX40 U9 ( .A(n8), .Y(n5) );
endmodule


module add_11 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   n29, temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_,
         temp2_0_, temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_,
         temp1_0_, n23, n24, n25, n27, n30, n31, n32, n33, n34;

  add_11_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n34, temp1_2_, 
        temp1_1_, n33}), .B({in2[6:3], n30, in2[1:0]}), .SUM(out3) );
  add_11_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, n31, temp2_3_, temp2_2_, 
        n25, temp2_0_}), .B(in), .SUM({n29, out1[5:0]}) );
  add_11_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n34, temp1_2_, 
        temp1_1_, n33}), .B({in3[6:2], n27, in3[0]}), .SUM(out2) );
  add_11_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n34, temp1_2_, 
        temp1_1_, n33}), .B({temp2_6_, temp2_5_, n31, temp2_3_, temp2_2_, n25, 
        temp2_0_}), .SUM(out) );
  add_11_DW01_add_4 add_30 ( .A({in2[6:3], n30, in2[1:0]}), .B({in3[6:2], n27, 
        in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_11_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2 U1 ( .A(in2[2]), .Y(n23) );
  BUFX2 U2 ( .A(temp1_0_), .Y(n24) );
  BUFX2 U3 ( .A(temp2_1_), .Y(n25) );
  BUFX10 U4 ( .A(n29), .Y(out1[6]) );
  BUFX4TH U5 ( .A(in3[1]), .Y(n27) );
  CLKBUFX40 U6 ( .A(n23), .Y(n30) );
  CLKBUFX40 U13 ( .A(temp2_4_), .Y(n31) );
  CLKINVX40 U14 ( .A(n24), .Y(n32) );
  CLKINVX40 U15 ( .A(n32), .Y(n33) );
  CLKBUFX40 U16 ( .A(temp1_3_), .Y(n34) );
endmodule


module tc_sm_47 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n25, n27, n28, n29, n30, n31, n32;

  CLKBUFX4 U3 ( .A(in[6]), .Y(n25) );
  NOR3X1TH U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U5 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U6 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U7 ( .A(in[2]), .Y(n31) );
  XNOR2XLTH U8 ( .A(n31), .B(n11), .Y(n10) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U10 ( .A(n25), .Y(n27) );
  OAI33X4TH U11 ( .A0(in[4]), .A1(n25), .A2(in[5]), .B0(n13), .B1(n28), .B2(
        n29), .Y(n8) );
  INVXLTH U12 ( .A(in[5]), .Y(n28) );
  INVXLTH U13 ( .A(in[4]), .Y(n29) );
  CLKINVX1TH U14 ( .A(in[3]), .Y(n30) );
  CLKBUFX1TH U15 ( .A(n25), .Y(out[4]) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U17 ( .A0(n27), .A1(n12), .B0(n25), .B1(n32), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U18 ( .A0(n27), .A1(n10), .B0(n25), .B1(n31), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U19 ( .A0(n9), .A1(n30), .B0(n25), .Y(n7) );
  OAI211XLTH U20 ( .A0(n25), .A1(n30), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U21 ( .A0N(n30), .A1N(n9), .B0(n25), .Y(n13) );
endmodule


module tc_sm_46 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n33, n34, n35, n36, n37, n38;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OAI221X2 U3 ( .A0(n35), .A1(n8), .B0(in[6]), .B1(n37), .C0(n6), .Y(out[2])
         );
  NAND3XL U4 ( .A(n33), .B(n34), .C(n6), .Y(out[1]) );
  AOI2BB1X4 U5 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  INVX2 U6 ( .A(in[6]), .Y(n35) );
  OAI211XL U8 ( .A0(in[6]), .A1(n36), .B0(n5), .C0(n6), .Y(out[3]) );
  AOI21X6 U9 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n6) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U11 ( .A(in[6]), .Y(out[4]) );
  OR2XLTH U12 ( .A(in[6]), .B(n38), .Y(n34) );
  OR2XLTH U13 ( .A(n35), .B(n10), .Y(n33) );
  XOR2XLTH U14 ( .A(in[0]), .B(n38), .Y(n10) );
  INVXLTH U15 ( .A(in[2]), .Y(n37) );
  XOR2XLTH U16 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI21XLTH U18 ( .A0(n7), .A1(n36), .B0(in[6]), .Y(n5) );
  INVXLTH U19 ( .A(in[3]), .Y(n36) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  INVXLTH U21 ( .A(in[1]), .Y(n38) );
endmodule


module tc_sm_45 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n19, n21, n22, n23, n24, n25,
         n26;

  OA21XLTH U3 ( .A0(in[6]), .A1(n24), .B0(n7), .Y(n18) );
  NAND2X2 U4 ( .A(n18), .B(n19), .Y(out[3]) );
  BUFX5 U5 ( .A(n8), .Y(n19) );
  OAI2BB1X1TH U6 ( .A0N(n24), .A1N(n9), .B0(in[6]), .Y(n13) );
  NAND2BXL U7 ( .AN(in[0]), .B(n19), .Y(out[0]) );
  OAI221XL U8 ( .A0(n21), .A1(n12), .B0(in[6]), .B1(n26), .C0(n19), .Y(out[1])
         );
  OAI221XL U9 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n25), .C0(n19), .Y(out[2])
         );
  INVXLTH U10 ( .A(in[6]), .Y(n21) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n24) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U14 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U16 ( .A(n25), .B(n11), .Y(n10) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U18 ( .A(in[2]), .Y(n25) );
  OAI21XLTH U19 ( .A0(n9), .A1(n24), .B0(in[6]), .Y(n7) );
  INVX2 U20 ( .A(in[5]), .Y(n22) );
  OAI33X4 U21 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n22), .B2(
        n23), .Y(n8) );
  INVXL U22 ( .A(in[4]), .Y(n23) );
endmodule


module tc_sm_44 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n30, n32, n33, n34, n35;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  INVXLTH U3 ( .A(in[6]), .Y(n32) );
  AOI21BX4 U4 ( .A0(in[6]), .A1(n11), .B0N(n30), .Y(n6) );
  NOR3X1TH U5 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U6 ( .A(in[6]), .Y(out[4]) );
  XOR2XLTH U8 ( .A(in[0]), .B(n35), .Y(n10) );
  INVXLTH U9 ( .A(in[1]), .Y(n35) );
  INVXLTH U10 ( .A(in[2]), .Y(n34) );
  XOR2XLTH U11 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI211XLTH U13 ( .A0(in[6]), .A1(n33), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI21XLTH U14 ( .A0(n7), .A1(n33), .B0(in[6]), .Y(n5) );
  INVXLTH U15 ( .A(in[3]), .Y(n33) );
  OAI21BX1 U16 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n30) );
  OAI221XLTH U17 ( .A0(n32), .A1(n8), .B0(in[6]), .B1(n34), .C0(n6), .Y(out[2]) );
  OAI221XLTH U18 ( .A0(n32), .A1(n10), .B0(in[6]), .B1(n35), .C0(n6), .Y(
        out[1]) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n6), .Y(out[0]) );
endmodule


module total_3_test_36 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n54, w5_4_, n4, n41, n43, n44, n45, n46, n47, n48, n49, n50, n51;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_47 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_46 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_45 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_44 sm_tc_4 ( .out(in1), .in(in) );
  add_11 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_47 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_46 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_45 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_44 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n47), .CK(clk), .RN(n4), .Q(
        h) );
  SDFFRQX1 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up1[2]) );
  SDFFRQXL up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n43), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n46), .CK(clk), .RN(rst), .Q(
        up1[0]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(n54) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n46), .CK(clk), .RN(rst), 
        .Q(up1[4]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up2[4]) );
  SDFFRQXL up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up1[1]) );
  SDFFRQX2 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n45), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  SDFFRQX1 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n45), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRQX2 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up2[3]) );
  SDFFRQX2 up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQX2 up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  CLKBUFX4TH U3 ( .A(rst), .Y(n4) );
  SDFFRX4 up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up3[3]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n43), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  DLY1X1TH U36 ( .A(n44), .Y(n41) );
  DLY1X1TH U37 ( .A(n54), .Y(up3[0]) );
  INVXLTH U38 ( .A(n44), .Y(n43) );
  DLY1X1TH U39 ( .A(n48), .Y(n44) );
  INVXLTH U40 ( .A(n44), .Y(n45) );
  INVXLTH U41 ( .A(n48), .Y(n46) );
  DLY1X1TH U42 ( .A(test_se), .Y(n47) );
  INVXLTH U43 ( .A(test_se), .Y(n48) );
  INVXLTH U44 ( .A(n41), .Y(n49) );
  INVXLTH U45 ( .A(n41), .Y(n50) );
  INVXLTH U46 ( .A(n44), .Y(n51) );
endmodule


module sm_tc_43 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n21, n22, n26, n27, n30;

  BUFX10 U2 ( .A(in[4]), .Y(n21) );
  CLKBUFX2TH U3 ( .A(in[1]), .Y(n22) );
  INVX4TH U4 ( .A(n21), .Y(n26) );
  XNOR2X1 U5 ( .A(n27), .B(n8), .Y(n5) );
  NOR2X4 U6 ( .A(n22), .B(in[0]), .Y(n8) );
  CLKBUFX1TH U7 ( .A(out[4]), .Y(out[6]) );
  INVX2 U8 ( .A(in[2]), .Y(n27) );
  AO21X1TH U9 ( .A0(in[0]), .A1(n22), .B0(n8), .Y(n6) );
  OAI2BB2X1TH U10 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  OAI22X4 U13 ( .A0(n21), .A1(n27), .B0(n26), .B1(n5), .Y(out[2]) );
  AOI31X2TH U14 ( .A0(n3), .A1(n5), .A2(n4), .B0(n26), .Y(out[4]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[5]) );
  BUFX2TH U18 ( .A(in[0]), .Y(out[0]) );
  AO2B2X4 U11 ( .B0(n22), .B1(n26), .A0(n21), .A1N(n6), .Y(out[1]) );
  XOR2X1 U12 ( .A(n30), .B(in[3]), .Y(n4) );
  CLKAND2X12 U15 ( .A(n8), .B(n27), .Y(n30) );
endmodule


module sm_tc_42 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n25, n26, n27, n28, n32, n33, n36;

  CLKBUFX1TH U2 ( .A(out[4]), .Y(out[6]) );
  CLKNAND2X4 U3 ( .A(n27), .B(n28), .Y(n5) );
  XNOR2X2 U4 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X2 U5 ( .B0(n32), .B1(n6), .A0N(in[1]), .A1N(n32), .Y(out[1]) );
  INVX6 U6 ( .A(in[4]), .Y(n32) );
  OAI22XLTH U7 ( .A0(in[4]), .A1(n33), .B0(n32), .B1(n5), .Y(out[2]) );
  NOR2X4TH U8 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX2TH U9 ( .A(in[2]), .Y(n33) );
  CLKBUFX2TH U10 ( .A(in[0]), .Y(out[0]) );
  NOR2BXL U12 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U13 ( .A(n33), .Y(n25) );
  NAND2XLTH U14 ( .A(n33), .B(n8), .Y(n27) );
  INVXLTH U15 ( .A(n8), .Y(n26) );
  OAI2BB2X1TH U16 ( .B0(n32), .B1(n4), .A0N(in[3]), .A1N(n32), .Y(out[3]) );
  AOI31X4 U17 ( .A0(n3), .A1(n4), .A2(n5), .B0(n32), .Y(out[4]) );
  NAND2XLTH U18 ( .A(n8), .B(n33), .Y(n7) );
  CLKBUFX1TH U19 ( .A(out[4]), .Y(out[5]) );
  AO21XLTH U20 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  AND2X8 U11 ( .A(n25), .B(n26), .Y(n36) );
  CLKINVX40 U21 ( .A(n36), .Y(n28) );
endmodule


module sm_tc_41 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n22, n24, n25, n29, n30, n33, n34, n35, n36, n37,
         n38;

  OAI2BB2X1 U4 ( .B0(n34), .B1(n4), .A0N(in[3]), .A1N(n34), .Y(out[3]) );
  OAI22X1 U7 ( .A0(n36), .A1(n30), .B0(n34), .B1(n5), .Y(out[2]) );
  NAND2XLTH U8 ( .A(n30), .B(n8), .Y(n24) );
  AOI31X4 U9 ( .A0(n3), .A1(n4), .A2(n5), .B0(n34), .Y(out[4]) );
  INVX5 U11 ( .A(in[4]), .Y(n29) );
  NAND2X5 U12 ( .A(n24), .B(n25), .Y(n5) );
  CLKNAND2X2 U13 ( .A(n22), .B(n37), .Y(n25) );
  CLKBUFX2TH U14 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[6]) );
  INVX2 U16 ( .A(in[2]), .Y(n30) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U20 ( .A(n30), .Y(n22) );
  CLKBUFX1TH U21 ( .A(out[4]), .Y(out[5]) );
  CLKINVX40 U2 ( .A(n29), .Y(n33) );
  CLKINVX40 U3 ( .A(n33), .Y(n34) );
  AOI21BX4 U5 ( .A0(in[0]), .A1(in[1]), .B0N(n37), .Y(n35) );
  CLKINVX40 U6 ( .A(n35), .Y(n6) );
  CLKINVX40 U10 ( .A(n34), .Y(n36) );
  OR2X8 U18 ( .A(in[1]), .B(in[0]), .Y(n37) );
  CLKINVX40 U19 ( .A(n37), .Y(n8) );
  AO2B2X4 U22 ( .B0(in[1]), .B1(n34), .A0(n35), .A1N(n34), .Y(out[1]) );
  XOR2X1 U23 ( .A(n38), .B(in[3]), .Y(n4) );
  CLKAND2X12 U24 ( .A(n8), .B(n30), .Y(n38) );
endmodule


module sm_tc_40 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  AOI31X1 U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  XNOR2X1 U3 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX1TH U4 ( .A(in[0]), .Y(out[0]) );
  NOR2X2TH U5 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U6 ( .A(in[2]), .Y(n21) );
  XNOR2X1TH U7 ( .A(n21), .B(n8), .Y(n5) );
  CLKINVX2TH U8 ( .A(in[4]), .Y(n22) );
  NAND2XLTH U9 ( .A(n8), .B(n21), .Y(n7) );
  INVXLTH U10 ( .A(out[4]), .Y(n18) );
  OAI22X1TH U11 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  INVXLTH U12 ( .A(n18), .Y(out[5]) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2BB2X1TH U14 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  INVXLTH U15 ( .A(n18), .Y(out[6]) );
  OAI2BB2XL U16 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_10_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3;
  wire   [6:2] carry;

  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR3X2 U3 ( .A(n3), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
  CLKINVX40 U5 ( .A(A[6]), .Y(n3) );
endmodule


module add_10_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_10_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_10_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X2 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_10_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_10 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         add_30_n14, add_30_n13, add_30_n10, add_30_n9, add_30_n6, add_30_n5,
         add_30_n4, add_30_n3, add_30_n2, add_30_n1, add_30_carry_2_,
         add_30_carry_3_, add_30_carry_4_, add_30_carry_5_, add_30_carry_6_,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32;

  add_10_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in2[6:3], n24, n23, in2[0]}), 
        .SUM(out3) );
  add_10_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_10_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in3[6:3], n32, n25, in3[0]}), 
        .SUM(out2) );
  add_10_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, 
        temp2_3_, temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_10_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  INVX2 U1 ( .A(add_30_n5), .Y(n28) );
  NAND3X2 U2 ( .A(add_30_n2), .B(add_30_n3), .C(add_30_n4), .Y(add_30_carry_5_) );
  ADDFHX2 U3 ( .A(n23), .B(n25), .CI(add_30_n6), .CO(add_30_carry_2_), .S(
        temp2_1_) );
  BUFX3 U4 ( .A(in2[2]), .Y(n24) );
  NAND2X4TH U5 ( .A(add_30_n13), .B(add_30_n14), .Y(temp2_0_) );
  XOR2X1 U6 ( .A(in2[6]), .B(in3[6]), .Y(add_30_n5) );
  XOR2X1 U11 ( .A(add_30_n1), .B(add_30_carry_4_), .Y(temp2_4_) );
  BUFX6 U13 ( .A(in2[1]), .Y(n23) );
  BUFX2 U14 ( .A(in3[1]), .Y(n25) );
  ADDFHX4 U15 ( .A(in2[3]), .B(in3[3]), .CI(add_30_carry_3_), .CO(
        add_30_carry_4_), .S(temp2_3_) );
  NAND2XL U17 ( .A(n28), .B(add_30_carry_6_), .Y(add_30_n10) );
  ADDFHX4 U18 ( .A(in2[5]), .B(in3[5]), .CI(add_30_carry_5_), .CO(
        add_30_carry_6_), .S(temp2_5_) );
  NAND2XLTH U20 ( .A(in3[4]), .B(in2[4]), .Y(add_30_n4) );
  CLKNAND2X2 U21 ( .A(add_30_carry_4_), .B(in2[4]), .Y(add_30_n3) );
  XOR2XLTH U22 ( .A(in2[4]), .B(in3[4]), .Y(add_30_n1) );
  ADDFHX4 U23 ( .A(n24), .B(n32), .CI(add_30_carry_2_), .CO(add_30_carry_3_), 
        .S(temp2_2_) );
  INVXLTH U24 ( .A(in2[0]), .Y(n26) );
  INVXLTH U25 ( .A(add_30_carry_6_), .Y(n29) );
  AND2XLTH U26 ( .A(in3[0]), .B(in2[0]), .Y(add_30_n6) );
  NAND2XLTH U27 ( .A(n27), .B(in2[0]), .Y(add_30_n14) );
  NAND2XLTH U28 ( .A(in3[0]), .B(n26), .Y(add_30_n13) );
  INVXLTH U29 ( .A(in3[0]), .Y(n27) );
  NAND2X2 U30 ( .A(add_30_n5), .B(n29), .Y(add_30_n9) );
  AND2X8 U16 ( .A(add_30_n9), .B(add_30_n10), .Y(n30) );
  CLKINVX40 U19 ( .A(n30), .Y(temp2_6_) );
  AND2X8 U31 ( .A(add_30_carry_4_), .B(in3[4]), .Y(n31) );
  CLKINVX40 U32 ( .A(n31), .Y(add_30_n2) );
  CLKBUFX40 U33 ( .A(in3[2]), .Y(n32) );
endmodule


module tc_sm_43 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n28) );
  XNOR2XLTH U7 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(in[6]), .Y(n24) );
  INVXLTH U10 ( .A(in[5]), .Y(n25) );
  INVXLTH U11 ( .A(in[4]), .Y(n26) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n27) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  OAI33X4TH U14 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U16 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_42 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n8, n9, n10, n11, n12, n13, n23, n24, n25, n27, n28, n29, n30, n31,
         n32, n33, n35, n36;

  OAI31X4 U3 ( .A0(n33), .A1(in[3]), .A2(in[2]), .B0(in[6]), .Y(n13) );
  OAI221X1 U4 ( .A0(n27), .A1(n8), .B0(in[6]), .B1(n30), .C0(n25), .Y(out[3])
         );
  CLKINVX1 U5 ( .A(in[6]), .Y(n27) );
  INVXLTH U7 ( .A(in[0]), .Y(n23) );
  CLKINVX1TH U8 ( .A(n23), .Y(n24) );
  OAI33X4 U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n29), .B2(n28), .Y(n9) );
  OAI221XL U10 ( .A0(n27), .A1(n11), .B0(in[6]), .B1(n31), .C0(n25), .Y(out[2]) );
  BUFX10 U11 ( .A(n9), .Y(n25) );
  INVXLTH U12 ( .A(n10), .Y(n33) );
  NOR2X1TH U13 ( .A(in[1]), .B(n24), .Y(n10) );
  CLKINVX1TH U14 ( .A(in[2]), .Y(n31) );
  INVXLTH U15 ( .A(in[4]), .Y(n29) );
  INVXLTH U16 ( .A(in[5]), .Y(n28) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U18 ( .AN(n24), .B(n25), .Y(out[0]) );
  INVXLTH U19 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U20 ( .A(n24), .B(in[1]), .Y(n12) );
  XNOR2XLTH U21 ( .A(n31), .B(n10), .Y(n11) );
  AOI21XLTH U22 ( .A0(n10), .A1(n31), .B0(n30), .Y(n8) );
  INVXLTH U23 ( .A(in[3]), .Y(n30) );
  OR2X8 U6 ( .A(n27), .B(n12), .Y(n35) );
  OR2X8 U24 ( .A(in[6]), .B(n32), .Y(n36) );
  NAND3X8 U25 ( .A(n35), .B(n36), .C(n25), .Y(out[1]) );
endmodule


module tc_sm_41 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n20, n21, n22, n23, n24, n25;

  BUFX10 U3 ( .A(n8), .Y(n18) );
  OAI2BB1X2 U4 ( .A0N(n23), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI211X2TH U5 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n18), .Y(out[3]) );
  OAI221X2 U6 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n18), .Y(out[2])
         );
  NAND2BX1 U7 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  OAI221X2 U8 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n18), .Y(out[1])
         );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U11 ( .A(in[4]), .Y(n22) );
  INVX1TH U12 ( .A(in[5]), .Y(n21) );
  INVXLTH U13 ( .A(in[6]), .Y(n20) );
  XNOR2XLTH U14 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[2]), .Y(n24) );
  OAI21XLTH U17 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  INVXLTH U18 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  CLKBUFX1TH U20 ( .A(in[6]), .Y(out[4]) );
  OAI33X4 U21 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n21), .B2(
        n22), .Y(n8) );
endmodule


module tc_sm_40 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n26, n27, n28, n29, n31;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  INVX1TH U3 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U4 ( .A0(n26), .A1(n8), .B0(in[6]), .B1(n28), .C0(n6), .Y(out[2])
         );
  NOR3X1TH U5 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  INVXLTH U6 ( .A(in[2]), .Y(n28) );
  XOR2XLTH U8 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n9) );
  XOR2XLTH U11 ( .A(in[0]), .B(n29), .Y(n10) );
  INVXLTH U12 ( .A(in[1]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  AOI21X8 U14 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n6) );
  AOI2BB1X4 U15 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  OAI221XLTH U16 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n29), .C0(n6), .Y(
        out[1]) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  OAI211XLTH U18 ( .A0(in[6]), .A1(n27), .B0(n5), .C0(n6), .Y(out[3]) );
  INVXLTH U19 ( .A(in[3]), .Y(n27) );
  OA21X4 U10 ( .A0(n7), .A1(n27), .B0(in[6]), .Y(n31) );
  CLKINVX40 U20 ( .A(n31), .Y(n5) );
endmodule


module total_3_test_37 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n56, n57, w5_4_, n4, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n52;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_43 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_42 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_41 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_40 sm_tc_4 ( .out(in1), .in(in) );
  add_10 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), 
        .in2(b1), .in3(c1), .in(in1) );
  tc_sm_43 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_42 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_41 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_40 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n45), .CK(clk), .RN(n4), 
        .Q(n57) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n44), .CK(clk), .RN(n4), .Q(
        h) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n40), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n41), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n47), .CK(clk), .RN(n4), .Q(
        up1[0]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n40), .CK(clk), .RN(n4), 
        .Q(n56) );
  SDFFRQX1TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up2[4]) );
  SDFFRQXLTH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n48), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n41), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n45), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRQX1TH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n48), .CK(clk), .RN(rst), 
        .Q(up1[1]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  SDFFRQX2 up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n44), .CK(clk), .RN(n4), 
        .Q(up1[4]) );
  CLKBUFX4TH U3 ( .A(rst), .Y(n4) );
  SDFFRHQX8 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n49), .CK(clk), .RN(rst), 
        .Q(n39) );
  INVXLTH U36 ( .A(n43), .Y(n40) );
  INVXLTH U37 ( .A(n42), .Y(n41) );
  DLY1X1TH U38 ( .A(n46), .Y(n42) );
  DLY1X1TH U39 ( .A(n46), .Y(n43) );
  INVXLTH U40 ( .A(n43), .Y(n44) );
  INVXLTH U41 ( .A(n42), .Y(n45) );
  INVXLTH U42 ( .A(test_se), .Y(n46) );
  INVXLTH U43 ( .A(n43), .Y(n47) );
  INVXLTH U44 ( .A(n42), .Y(n48) );
  INVXLTH U45 ( .A(n43), .Y(n49) );
  INVXLTH U46 ( .A(n42), .Y(n50) );
  CLKINVX40 U47 ( .A(n39), .Y(n52) );
  CLKINVX40 U48 ( .A(n52), .Y(up1[2]) );
  DLY1X1TH U49 ( .A(n56), .Y(up2[3]) );
  DLY1X1TH U50 ( .A(n57), .Y(up3[3]) );
endmodule


module sm_tc_39 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n23;

  XNOR2X1 U2 ( .A(n23), .B(n8), .Y(n5) );
  NOR2X3 U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  AOI31X1 U4 ( .A0(n5), .A1(n4), .A2(n3), .B0(n22), .Y(out[4]) );
  XNOR2X2 U5 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X4 U6 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  OAI22X1 U7 ( .A0(in[4]), .A1(n23), .B0(n22), .B1(n5), .Y(out[2]) );
  INVX2TH U8 ( .A(in[2]), .Y(n23) );
  CLKINVX2TH U9 ( .A(in[4]), .Y(n22) );
  CLKBUFX1TH U10 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[6]) );
  NAND2XLTH U13 ( .A(n8), .B(n23), .Y(n7) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2BB2XLTH U15 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  AO21XLTH U16 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module sm_tc_38 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n4, n5, n6, n7, n8, n9, n20, n21, n23, n26, n27, n28, n31;

  NOR2XLTH U2 ( .A(in[4]), .B(n27), .Y(n20) );
  NOR2X2 U3 ( .A(n26), .B(n7), .Y(n21) );
  OR2X2 U4 ( .A(n20), .B(n21), .Y(out[2]) );
  INVX4 U5 ( .A(in[2]), .Y(n27) );
  INVX4 U6 ( .A(in[4]), .Y(n26) );
  AOI31X4 U8 ( .A0(n4), .A1(n28), .A2(n5), .B0(n26), .Y(out[4]) );
  OAI2B2X4 U9 ( .A1N(in[1]), .A0(in[4]), .B0(n6), .B1(n26), .Y(out[1]) );
  XOR2X1TH U10 ( .A(in[2]), .B(n9), .Y(n7) );
  XNOR2X1TH U11 ( .A(n8), .B(in[3]), .Y(n5) );
  AND2XLTH U12 ( .A(n6), .B(n7), .Y(n4) );
  XOR2X2TH U14 ( .A(in[1]), .B(n28), .Y(n6) );
  CLKBUFX1TH U15 ( .A(in[0]), .Y(out[0]) );
  INVX1TH U16 ( .A(out[4]), .Y(n23) );
  INVXLTH U17 ( .A(n23), .Y(out[6]) );
  INVXLTH U18 ( .A(in[0]), .Y(n28) );
  INVXLTH U19 ( .A(n23), .Y(out[5]) );
  NAND2XLTH U20 ( .A(n9), .B(n27), .Y(n8) );
  OR2X8 U7 ( .A(in[1]), .B(in[0]), .Y(n31) );
  CLKINVX40 U13 ( .A(n31), .Y(n9) );
  AO2B2X4 U21 ( .B0(in[3]), .B1(n26), .A0(in[4]), .A1N(n5), .Y(out[3]) );
endmodule


module sm_tc_37 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n4, n5, n6, n7, n8, n9, n21, n25, n26;

  OAI2BB2X2 U2 ( .B0(n25), .B1(n5), .A0N(in[3]), .A1N(n25), .Y(out[3]) );
  INVX4 U3 ( .A(n21), .Y(n25) );
  AO21X2 U4 ( .A0(in[0]), .A1(in[1]), .B0(n9), .Y(n7) );
  BUFX2 U5 ( .A(in[0]), .Y(out[0]) );
  NOR2X6 U6 ( .A(in[1]), .B(in[0]), .Y(n9) );
  XNOR2X2 U7 ( .A(n8), .B(in[3]), .Y(n5) );
  BUFX2 U8 ( .A(in[4]), .Y(n21) );
  OAI22X1 U9 ( .A0(n21), .A1(n26), .B0(n6), .B1(n25), .Y(out[2]) );
  NAND2X1TH U10 ( .A(n9), .B(n26), .Y(n8) );
  OAI2BB2X2 U11 ( .B0(n25), .B1(n7), .A0N(in[1]), .A1N(n25), .Y(out[1]) );
  AOI31X2TH U12 ( .A0(n4), .A1(n5), .A2(n6), .B0(n25), .Y(out[4]) );
  CLKINVX1TH U13 ( .A(in[2]), .Y(n26) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[6]) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U17 ( .AN(n7), .B(in[0]), .Y(n4) );
  XOR2X1 U15 ( .A(in[2]), .B(n9), .Y(n6) );
endmodule


module sm_tc_36 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  NAND2X1TH U2 ( .A(n8), .B(n21), .Y(n7) );
  CLKBUFX1TH U3 ( .A(in[0]), .Y(out[0]) );
  AOI31X4TH U4 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  XNOR2X2TH U5 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKINVX2TH U6 ( .A(in[4]), .Y(n22) );
  OAI2BB2X2TH U7 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  INVXLTH U8 ( .A(n18), .Y(out[6]) );
  OAI22X2TH U9 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  NOR2X1TH U10 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n21) );
  OAI2BB2X1TH U12 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  INVXLTH U13 ( .A(out[4]), .Y(n18) );
  INVXLTH U14 ( .A(n18), .Y(out[5]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  XNOR2X1TH U16 ( .A(n21), .B(n8), .Y(n5) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_9_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X8 U3 ( .A(n4), .B(A[6]), .Y(n2) );
  CLKXOR2X8 U4 ( .A(n2), .B(carry[6]), .Y(n3) );
  CLKINVX40 U5 ( .A(n3), .Y(SUM[6]) );
  CLKINVX40 U6 ( .A(B[6]), .Y(n4) );
endmodule


module add_9_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHX2TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_9_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X2 U3 ( .A(B[6]), .B(A[6]), .Y(n2) );
  CLKXOR2X12 U4 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
endmodule


module add_9_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n3;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR2X4TH U2 ( .A(n3), .B(carry[6]), .Y(SUM[6]) );
  XNOR2XLTH U3 ( .A(A[6]), .B(B[6]), .Y(n3) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_9_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3XL U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_9_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n4, n5, n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1TH U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(n5) );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(n4) );
  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKBUFX40 U3 ( .A(n4), .Y(SUM[5]) );
  CLKBUFX40 U4 ( .A(n5), .Y(SUM[4]) );
endmodule


module add_9 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n22, n23, n24, n25, n26, n27;

  add_9_DW01_add_0 add_34 ( .A({n25, temp1_5_, temp1_4_, n26, temp1_2_, 
        temp1_1_, temp1_0_}), .B({n27, in2[5:2], n23, n22}), .SUM(out3) );
  add_9_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_9_DW01_add_2 add_32 ( .A({n25, temp1_5_, temp1_4_, n26, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in3[6:2], n24, in3[0]}), .SUM(out2) );
  add_9_DW01_add_3 add_31 ( .A({n25, temp1_5_, temp1_4_, n26, temp1_2_, 
        temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_9_DW01_add_4 add_30 ( .A({n27, in2[5:2], n23, in2[0]}), .B(in3), .SUM({
        temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_})
         );
  add_9_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2 U1 ( .A(in2[0]), .Y(n22) );
  CLKBUFX2 U2 ( .A(in2[1]), .Y(n23) );
  CLKBUFX2TH U3 ( .A(in3[1]), .Y(n24) );
  CLKBUFX40 U4 ( .A(temp1_6_), .Y(n25) );
  CLKBUFX40 U5 ( .A(temp1_3_), .Y(n26) );
  CLKBUFX40 U6 ( .A(in2[6]), .Y(n27) );
endmodule


module tc_sm_39 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n27, n28, n29, n30, n31, n32;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n31) );
  XNOR2XLTH U7 ( .A(n31), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(in[6]), .Y(n27) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n28), .B2(
        n29), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n29) );
  INVXLTH U12 ( .A(in[5]), .Y(n28) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n30) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI21XLTH U16 ( .A0(n9), .A1(n30), .B0(in[6]), .Y(n7) );
  OAI221XLTH U17 ( .A0(n27), .A1(n12), .B0(in[6]), .B1(n32), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U18 ( .A0(n27), .A1(n10), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[2]) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n30), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n30), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_38 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n19, n20, n21, n23, n24, n25, n26,
         n27, n28;

  BUFX10 U3 ( .A(n8), .Y(n19) );
  OAI2BB1X1 U4 ( .A0N(n26), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI211XLTH U5 ( .A0(in[6]), .A1(n26), .B0(n7), .C0(n19), .Y(out[3]) );
  OR2XLTH U6 ( .A(n23), .B(n12), .Y(n20) );
  OR2XLTH U7 ( .A(in[6]), .B(n28), .Y(n21) );
  NAND3XL U8 ( .A(n20), .B(n21), .C(n19), .Y(out[1]) );
  OAI221X2TH U9 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n27), .C0(n19), .Y(
        out[2]) );
  NAND2BX1TH U10 ( .AN(in[0]), .B(n19), .Y(out[0]) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n26) );
  INVXLTH U12 ( .A(in[4]), .Y(n25) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U15 ( .A(n27), .B(n11), .Y(n10) );
  OAI21XLTH U16 ( .A0(n9), .A1(n26), .B0(in[6]), .Y(n7) );
  INVX2 U17 ( .A(in[5]), .Y(n24) );
  INVXLTH U18 ( .A(in[6]), .Y(n23) );
  INVXLTH U19 ( .A(in[1]), .Y(n28) );
  XNOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U22 ( .A(in[2]), .Y(n27) );
  OAI33X4 U23 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n24), .B2(
        n25), .Y(n8) );
endmodule


module tc_sm_37 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n26, n27,
         n28;

  OAI211XL U4 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221XL U5 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1])
         );
  OAI221XL U6 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2])
         );
  INVX2TH U7 ( .A(in[4]), .Y(n21) );
  INVX1TH U8 ( .A(in[5]), .Y(n20) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n22) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U11 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U12 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U14 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[2]), .Y(n23) );
  OAI21XLTH U17 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  INVXLTH U18 ( .A(in[6]), .Y(n19) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  AOI33X4 U3 ( .A0(n21), .A1(n27), .A2(n20), .B0(n28), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U20 ( .A(n26), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n27) );
  AOI21BX4 U22 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n28) );
endmodule


module tc_sm_36 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n19, n21, n22, n23, n24, n26, n27, n28;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OAI221XL U3 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n24), .C0(n6), .Y(out[1])
         );
  CLKINVX2 U4 ( .A(in[6]), .Y(n21) );
  AOI21BX4 U5 ( .A0(in[6]), .A1(n11), .B0N(n19), .Y(n6) );
  OAI21BX4 U6 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n19) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U9 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U10 ( .A0(n7), .A1(n22), .B0(in[6]), .Y(n5) );
  INVXLTH U11 ( .A(in[3]), .Y(n22) );
  XOR2XLTH U12 ( .A(in[0]), .B(n24), .Y(n10) );
  INVXLTH U13 ( .A(in[1]), .Y(n24) );
  INVXLTH U14 ( .A(in[2]), .Y(n23) );
  XOR2XLTH U15 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n9) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  OR2X8 U17 ( .A(n21), .B(n8), .Y(n26) );
  OR2X8 U19 ( .A(in[6]), .B(n23), .Y(n27) );
  NAND3X8 U20 ( .A(n26), .B(n27), .C(n6), .Y(out[2]) );
  OAI2B11X4 U21 ( .A1N(n28), .A0(n22), .B0(n5), .C0(n6), .Y(out[3]) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n28) );
endmodule


module total_3_test_38 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n4, n39, n40, n41, n42, n43, n44, n45, n46, n47;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_39 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_38 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_37 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_36 sm_tc_4 ( .out(in1), .in(in) );
  add_9 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), .in2(
        b1), .in3(c1), .in(in1) );
  tc_sm_39 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_38 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_37 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_36 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n41), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n40), .CK(clk), .RN(n4), .Q(
        h) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n42), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRQX1TH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRQX2TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n43), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n46), .CK(clk), .RN(n4), .Q(
        up1[0]) );
  SDFFRQX1TH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n43), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  SDFFRHQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n42), .CK(clk), .RN(n44), .Q(up1[4]) );
  SDFFRHQX1TH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n43), .CK(clk), .RN(n44), .Q(up3[3]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n42), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRHQX1TH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n46), .CK(clk), .RN(n4), 
        .Q(up1[1]) );
  SDFFRHQX1TH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n47), .CK(clk), .RN(n4), 
        .Q(up2[3]) );
  SDFFRQX4 up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n41), .CK(clk), .RN(rst), 
        .Q(up2[4]) );
  CLKBUFX4TH U3 ( .A(rst), .Y(n4) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n42), .CK(clk), .RN(n4), 
        .Q(up1[2]) );
  SDFFRHQX8 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n43), .CK(clk), .RN(n4), 
        .Q(up1[3]) );
  SDFFRX4 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n40), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  DLY1X1TH U36 ( .A(n45), .Y(n39) );
  INVXLTH U37 ( .A(n39), .Y(n40) );
  INVXLTH U38 ( .A(n39), .Y(n41) );
  DLY1X1TH U39 ( .A(test_se), .Y(n42) );
  DLY1X1TH U40 ( .A(test_se), .Y(n43) );
  DLY1X1TH U41 ( .A(n4), .Y(n44) );
  INVXLTH U42 ( .A(test_se), .Y(n45) );
  INVXLTH U43 ( .A(n39), .Y(n46) );
  INVXLTH U44 ( .A(n39), .Y(n47) );
endmodule


module sm_tc_35 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n22, n27, n30, n31, n32, n33;

  CLKBUFX2TH U2 ( .A(in[0]), .Y(out[0]) );
  BUFX2TH U3 ( .A(in[4]), .Y(n22) );
  AOI31X1 U6 ( .A0(n3), .A1(n4), .A2(n5), .B0(n33), .Y(out[4]) );
  CLKBUFX1TH U7 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X4 U9 ( .B0(n33), .B1(n6), .A0N(in[1]), .A1N(n33), .Y(out[1]) );
  NOR2X6 U10 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX2TH U11 ( .A(in[2]), .Y(n27) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2XLTH U13 ( .B0(n33), .B1(n4), .A0N(in[3]), .A1N(n33), .Y(out[3]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2B2X2 U4 ( .A1N(n31), .A0(n5), .B0(n31), .B1(n27), .Y(out[2]) );
  XNOR2X1 U5 ( .A(n27), .B(n8), .Y(n5) );
  CLKINVX40 U8 ( .A(n22), .Y(n30) );
  CLKINVX40 U14 ( .A(n30), .Y(n31) );
  XOR2X1 U16 ( .A(n32), .B(in[3]), .Y(n4) );
  CLKAND2X12 U18 ( .A(n8), .B(n27), .Y(n32) );
  CLKINVX40 U19 ( .A(n31), .Y(n33) );
endmodule


module sm_tc_34 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n24, n28, n29, n32, n33, n34, n35, n36;

  BUFX2 U2 ( .A(in[4]), .Y(n24) );
  OAI2BB2X2 U3 ( .B0(n36), .B1(n6), .A0N(in[1]), .A1N(n36), .Y(out[1]) );
  BUFX2 U5 ( .A(n34), .Y(out[0]) );
  INVX2 U6 ( .A(n24), .Y(n28) );
  OAI2BB2X2TH U8 ( .B0(n36), .B1(n4), .A0N(in[3]), .A1N(n36), .Y(out[3]) );
  INVX1TH U9 ( .A(in[2]), .Y(n29) );
  CLKBUFX1TH U10 ( .A(out[4]), .Y(out[6]) );
  AO21X1TH U12 ( .A0(n34), .A1(in[1]), .B0(n8), .Y(n6) );
  AOI31X2TH U14 ( .A0(n3), .A1(n4), .A2(n5), .B0(n36), .Y(out[4]) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U16 ( .AN(n6), .B(n34), .Y(n3) );
  XNOR2X1TH U17 ( .A(n29), .B(n8), .Y(n5) );
  OR2X8 U4 ( .A(in[1]), .B(n34), .Y(n32) );
  CLKINVX40 U7 ( .A(n32), .Y(n8) );
  XNOR2X1 U11 ( .A(n33), .B(in[3]), .Y(n4) );
  CLKNAND2X12 U13 ( .A(n8), .B(n29), .Y(n33) );
  CLKBUFX40 U18 ( .A(in[0]), .Y(n34) );
  CLKINVX40 U19 ( .A(n28), .Y(n35) );
  CLKINVX40 U20 ( .A(n35), .Y(n36) );
  OAI2B2X4 U21 ( .A1N(n36), .A0(n29), .B0(n36), .B1(n5), .Y(out[2]) );
endmodule


module sm_tc_33 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n28, n29, n30, n31, n42, n35, n36, n39, n41;

  OAI2BB2X4 U2 ( .B0(n35), .B1(n6), .A0N(in[1]), .A1N(n35), .Y(out[1]) );
  BUFX2 U3 ( .A(in[4]), .Y(n31) );
  CLKBUFX1 U4 ( .A(out[4]), .Y(out[5]) );
  CLKNAND2X2TH U5 ( .A(n29), .B(n30), .Y(n4) );
  NAND2X2 U6 ( .A(n41), .B(n28), .Y(n30) );
  CLKBUFX2TH U7 ( .A(out[4]), .Y(out[6]) );
  INVX2TH U8 ( .A(n31), .Y(n35) );
  CLKBUFX2 U9 ( .A(in[0]), .Y(n42) );
  CLKNAND2X2TH U10 ( .A(n7), .B(in[3]), .Y(n29) );
  OAI2BB2X4TH U12 ( .B0(n35), .B1(n4), .A0N(in[3]), .A1N(n35), .Y(out[3]) );
  OAI22X1 U13 ( .A0(n31), .A1(n36), .B0(n35), .B1(n5), .Y(out[2]) );
  NOR2X8 U14 ( .A(in[1]), .B(out[0]), .Y(n8) );
  INVXLTH U15 ( .A(in[3]), .Y(n28) );
  AOI31X2 U16 ( .A0(n3), .A1(n4), .A2(n5), .B0(n35), .Y(out[4]) );
  CLKINVX1TH U18 ( .A(in[2]), .Y(n36) );
  AO21XLTH U20 ( .A0(out[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2BXLTH U21 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKINVX40 U11 ( .A(n42), .Y(n39) );
  CLKINVX40 U17 ( .A(n39), .Y(out[0]) );
  XOR2X1 U19 ( .A(in[2]), .B(n8), .Y(n5) );
  AND2X8 U22 ( .A(n8), .B(n36), .Y(n41) );
  CLKINVX40 U23 ( .A(n41), .Y(n7) );
endmodule


module sm_tc_32 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  AOI31X1 U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  INVX2 U3 ( .A(out[4]), .Y(n18) );
  NOR2X2TH U4 ( .A(in[1]), .B(in[0]), .Y(n8) );
  NAND2XLTH U5 ( .A(n8), .B(n21), .Y(n7) );
  CLKBUFX1TH U6 ( .A(in[0]), .Y(out[0]) );
  OAI22X1TH U7 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  INVXLTH U8 ( .A(n18), .Y(out[6]) );
  CLKINVX1TH U9 ( .A(in[2]), .Y(n21) );
  CLKINVX2TH U10 ( .A(in[4]), .Y(n22) );
  OAI2BB2X1TH U11 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  NOR2BXLTH U12 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U13 ( .A(n18), .Y(out[5]) );
  OAI2BB2X2TH U14 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  XNOR2X1TH U15 ( .A(n21), .B(n8), .Y(n5) );
  XNOR2X1TH U16 ( .A(n7), .B(in[3]), .Y(n4) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_8_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_8_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [6:2] carry;

  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2XLTH U2 ( .A(A[1]), .B(n1), .Y(n3) );
  NAND2XLTH U3 ( .A(n1), .B(B[1]), .Y(n5) );
  NAND3X2TH U4 ( .A(n5), .B(n4), .C(n3), .Y(carry[2]) );
  CLKXOR2X1TH U5 ( .A(n2), .B(A[1]), .Y(SUM[1]) );
  XOR2XLTH U6 ( .A(B[1]), .B(n1), .Y(n2) );
  NAND2XLTH U7 ( .A(A[1]), .B(B[1]), .Y(n4) );
  AND2X1TH U8 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U9 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n6) );
  CLKINVX40 U10 ( .A(n6), .Y(SUM[6]) );
endmodule


module add_8_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_8_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(B[1]), .B(A[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_8_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3XL U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  NAND3X2 U1 ( .A(n2), .B(n3), .C(n4), .Y(carry[4]) );
  NAND2X1 U3 ( .A(A[3]), .B(B[3]), .Y(n3) );
  NAND2XLTH U4 ( .A(A[3]), .B(carry[3]), .Y(n2) );
  XOR2XL U5 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U6 ( .A(carry[3]), .B(B[3]), .Y(n4) );
  AND2XLTH U7 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U2 ( .A(n5), .B(carry[3]), .C(B[3]), .Y(SUM[3]) );
  CLKINVX40 U8 ( .A(A[3]), .Y(n5) );
endmodule


module add_8_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_8 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n25, n26, n29, n30, n31, n32, n33, n34, n35;

  add_8_DW01_add_0 add_34 ( .A({temp1_6_, n33, temp1_4_, temp1_3_, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in2[6:4], n31, in2[2], n25, in2[0]}), .SUM(
        out3) );
  add_8_DW01_add_1 add_33 ( .A({temp2_6_, n30, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, n35}), .B(in), .SUM(out1) );
  add_8_DW01_add_2 add_32 ( .A({temp1_6_, n33, temp1_4_, temp1_3_, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in3[6:3], n26, n29, in3[0]}), .SUM(out2) );
  add_8_DW01_add_3 add_31 ( .A({temp1_6_, n33, temp1_4_, temp1_3_, temp1_2_, 
        temp1_1_, temp1_0_}), .B({temp2_6_, n30, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, n35}), .SUM(out) );
  add_8_DW01_add_4 add_30 ( .A({in2[6:4], n31, in2[2:0]}), .B({in3[6:3], n26, 
        n29, in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_8_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2TH U1 ( .A(in2[1]), .Y(n25) );
  BUFX2TH U2 ( .A(in3[2]), .Y(n26) );
  CLKBUFX2TH U3 ( .A(in3[1]), .Y(n29) );
  CLKBUFX40 U4 ( .A(temp2_5_), .Y(n30) );
  CLKBUFX40 U5 ( .A(in2[3]), .Y(n31) );
  CLKBUFX40 U6 ( .A(temp2_0_), .Y(n32) );
  CLKBUFX40 U13 ( .A(temp1_5_), .Y(n33) );
  CLKINVX40 U14 ( .A(n32), .Y(n34) );
  CLKINVX40 U15 ( .A(n34), .Y(n35) );
endmodule


module tc_sm_35 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U10 ( .A(in[4]), .Y(n28) );
  INVXLTH U11 ( .A(in[5]), .Y(n27) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_34 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n22, n23, n25, n26, n27, n28, n29,
         n30, n32, n33, n34;

  BUFX10 U3 ( .A(n8), .Y(n23) );
  OAI2BB1X4 U5 ( .A0N(n28), .A1N(n9), .B0(in[6]), .Y(n13) );
  OA21XL U6 ( .A0(in[6]), .A1(n28), .B0(n7), .Y(n22) );
  OAI221X1 U7 ( .A0(n25), .A1(n10), .B0(in[6]), .B1(n29), .C0(n23), .Y(out[2])
         );
  INVXLTH U8 ( .A(in[6]), .Y(n25) );
  OAI221X2 U9 ( .A0(n34), .A1(n12), .B0(in[6]), .B1(n30), .C0(n23), .Y(out[1])
         );
  NAND2XLTH U10 ( .A(n22), .B(n23), .Y(out[3]) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n28) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U14 ( .A(n29), .B(n11), .Y(n10) );
  INVXLTH U15 ( .A(in[2]), .Y(n29) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n23), .Y(out[0]) );
  INVX2 U17 ( .A(in[5]), .Y(n26) );
  INVXLTH U18 ( .A(in[1]), .Y(n30) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4 U21 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n26), .B2(
        n27), .Y(n8) );
  INVXL U22 ( .A(in[4]), .Y(n27) );
  AOI2BB1X4 U4 ( .A0N(n9), .A1N(n28), .B0(n33), .Y(n32) );
  CLKINVX40 U23 ( .A(n32), .Y(n7) );
  CLKINVX40 U24 ( .A(in[6]), .Y(n33) );
  INVXLTH U25 ( .A(in[6]), .Y(n34) );
endmodule


module tc_sm_33 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n21, n23, n24, n25, n26, n27,
         n28;

  AOI21BX2 U3 ( .A0(n26), .A1(n9), .B0N(in[6]), .Y(n21) );
  CLKINVX4TH U4 ( .A(n19), .Y(n8) );
  INVXLTH U5 ( .A(in[6]), .Y(n20) );
  AOI33X4 U6 ( .A0(n25), .A1(n20), .A2(n24), .B0(n21), .B1(in[5]), .B2(in[4]), 
        .Y(n19) );
  INVXLTH U7 ( .A(in[4]), .Y(n25) );
  INVXLTH U8 ( .A(in[5]), .Y(n24) );
  OAI211XL U9 ( .A0(in[6]), .A1(n26), .B0(n7), .C0(n8), .Y(out[3]) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n26) );
  INVXLTH U12 ( .A(in[6]), .Y(n23) );
  XNOR2XLTH U13 ( .A(n27), .B(n11), .Y(n10) );
  OAI21XLTH U14 ( .A0(n9), .A1(n26), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U17 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n27), .C0(n8), .Y(
        out[2]) );
  NOR2XLTH U18 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U19 ( .A(in[2]), .Y(n27) );
  OAI221XLTH U20 ( .A0(n23), .A1(n12), .B0(in[6]), .B1(n28), .C0(n8), .Y(
        out[1]) );
  INVXLTH U21 ( .A(in[1]), .Y(n28) );
  XNOR2XLTH U22 ( .A(in[0]), .B(in[1]), .Y(n12) );
endmodule


module tc_sm_32 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n22, n23, n24, n25, n27, n28, n29;

  OAI2B11X2TH U4 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  INVXLTH U5 ( .A(in[6]), .Y(n22) );
  OAI211XLTH U6 ( .A0(in[6]), .A1(n23), .B0(n5), .C0(n29), .Y(out[3]) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  INVXLTH U9 ( .A(in[2]), .Y(n24) );
  XOR2XLTH U10 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI21XLTH U12 ( .A0(n7), .A1(n23), .B0(in[6]), .Y(n5) );
  INVXLTH U13 ( .A(in[3]), .Y(n23) );
  XOR2XLTH U14 ( .A(in[0]), .B(n25), .Y(n10) );
  INVXLTH U15 ( .A(in[1]), .Y(n25) );
  CLKBUFX1TH U16 ( .A(in[6]), .Y(out[4]) );
  OAI221XLTH U17 ( .A0(n22), .A1(n8), .B0(in[6]), .B1(n24), .C0(n29), .Y(
        out[2]) );
  OAI221XLTH U18 ( .A0(n22), .A1(n10), .B0(in[6]), .B1(n25), .C0(n29), .Y(
        out[1]) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n29), .Y(out[0]) );
  AOI21BX4 U3 ( .A0(in[6]), .A1(n11), .B0N(n27), .Y(n6) );
  OAI21BX4 U7 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n27) );
  CLKINVX40 U20 ( .A(n6), .Y(n28) );
  CLKINVX40 U21 ( .A(n28), .Y(n29) );
endmodule


module total_3_test_39 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n4, n39, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52
;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_35 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_34 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_33 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_32 sm_tc_4 ( .out(in1), .in(in) );
  add_8 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), .in2(
        {b1[6], n39, b1[4:0]}), .in3(c1), .in(in1) );
  tc_sm_35 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_34 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_33 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_32 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n46), .CK(clk), .RN(n4), 
        .Q(up2[4]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up2[0]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n43), .CK(clk), .RN(rst), 
        .Q(h) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n46), .CK(clk), .RN(n4), 
        .Q(up3[3]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n47), .CK(clk), .RN(rst), 
        .Q(up1[3]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n51), .CK(clk), .RN(n4), 
        .Q(up2[3]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up3[2]) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n52), .CK(clk), .RN(n4), 
        .Q(up1[4]) );
  SDFFRQX2TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n42), .CK(clk), .RN(n4), 
        .Q(up3[4]) );
  SDFFRQX2TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n47), .CK(clk), .RN(n4), .Q(
        up1[0]) );
  SDFFRQX1TH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n43), .CK(clk), .RN(n4), 
        .Q(up1[1]) );
  SDFFRHQX2TH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up2[2]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up3[1]) );
  CLKBUFX4TH U3 ( .A(rst), .Y(n4) );
  SDFFRX4 up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n50), .CK(clk), .RN(n4), 
        .Q(up3[0]) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n49), .CK(clk), .RN(n4), 
        .Q(up2[1]) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n42), .CK(clk), .RN(n4), 
        .Q(up1[2]) );
  CLKBUFX40 U36 ( .A(b1[5]), .Y(n39) );
  INVXLTH U37 ( .A(n45), .Y(n42) );
  INVXLTH U38 ( .A(n44), .Y(n43) );
  DLY1X1TH U39 ( .A(n48), .Y(n44) );
  DLY1X1TH U40 ( .A(n48), .Y(n45) );
  INVXLTH U41 ( .A(n45), .Y(n46) );
  INVXLTH U42 ( .A(n44), .Y(n47) );
  INVXLTH U43 ( .A(test_se), .Y(n48) );
  INVXLTH U44 ( .A(n45), .Y(n49) );
  INVXLTH U45 ( .A(n44), .Y(n50) );
  INVXLTH U46 ( .A(n45), .Y(n51) );
  INVXLTH U47 ( .A(n44), .Y(n52) );
endmodule


module sm_tc_31 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n21, n25, n26, n29, n30, n31, n32, n33;

  AO21X2 U2 ( .A0(in[0]), .A1(n32), .B0(n8), .Y(n6) );
  NOR2X4 U3 ( .A(n32), .B(in[0]), .Y(n8) );
  OAI22X1 U5 ( .A0(n21), .A1(n25), .B0(n26), .B1(n5), .Y(out[2]) );
  AOI31X1 U6 ( .A0(n3), .A1(n29), .A2(n4), .B0(n26), .Y(out[4]) );
  INVX2TH U7 ( .A(in[2]), .Y(n25) );
  CLKBUFX2TH U9 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U10 ( .A(n26), .Y(n21) );
  INVX4TH U11 ( .A(in[4]), .Y(n26) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X2 U13 ( .B0(n26), .B1(n6), .A0N(n32), .A1N(n26), .Y(out[1]) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  XOR2X1 U4 ( .A(n25), .B(n30), .Y(n29) );
  XOR2X1 U8 ( .A(n25), .B(n30), .Y(n5) );
  CLKINVX40 U14 ( .A(n8), .Y(n30) );
  AO2B2BX4 U16 ( .A0(n31), .A1N(n4), .B0(in[3]), .B1N(n31), .Y(out[3]) );
  CLKINVX40 U18 ( .A(n26), .Y(n31) );
  CLKBUFX40 U19 ( .A(in[1]), .Y(n32) );
  XOR2X1 U20 ( .A(n33), .B(in[3]), .Y(n4) );
  CLKAND2X12 U21 ( .A(n8), .B(n25), .Y(n33) );
endmodule


module sm_tc_30 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n12, n13, n14, n15;

  AOI31X2 U2 ( .A0(n6), .A1(n3), .A2(n4), .B0(n12), .Y(out[4]) );
  XNOR2X1 U3 ( .A(n8), .B(in[3]), .Y(n3) );
  INVX2TH U5 ( .A(n14), .Y(n12) );
  OAI2BB2X4 U6 ( .B0(n12), .B1(n5), .A0N(in[1]), .A1N(n12), .Y(out[1]) );
  XNOR2X4TH U7 ( .A(n13), .B(n7), .Y(n4) );
  CLKBUFX1TH U8 ( .A(in[0]), .Y(out[0]) );
  CLKNAND2X4 U9 ( .A(n7), .B(n13), .Y(n8) );
  OAI2BB2X2TH U10 ( .B0(n12), .B1(n3), .A0N(in[3]), .A1N(n12), .Y(out[3]) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  OAI22X1TH U12 ( .A0(n14), .A1(n13), .B0(n12), .B1(n4), .Y(out[2]) );
  CLKINVX1TH U13 ( .A(in[2]), .Y(n13) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U15 ( .AN(n5), .B(in[0]), .Y(n6) );
  OAI2BB1X4 U4 ( .A0N(in[0]), .A1N(in[1]), .B0(n15), .Y(n5) );
  CLKBUFX40 U16 ( .A(in[4]), .Y(n14) );
  OR2X8 U17 ( .A(in[1]), .B(in[0]), .Y(n15) );
  CLKINVX40 U18 ( .A(n15), .Y(n7) );
endmodule


module sm_tc_29 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n38, n3, n4, n5, n6, n7, n8, n19, n20, n21, n22, n23, n27, n28, n30,
         n31, n32, n33, n34, n35, n37;

  INVX4 U2 ( .A(n27), .Y(n19) );
  NAND2XLTH U3 ( .A(n27), .B(n8), .Y(n21) );
  NAND2X4 U4 ( .A(n19), .B(n20), .Y(n22) );
  CLKNAND2X8 U5 ( .A(n21), .B(n22), .Y(n5) );
  INVXLTH U6 ( .A(n8), .Y(n20) );
  INVX4 U7 ( .A(in[2]), .Y(n27) );
  NOR2X6 U8 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI22XLTH U9 ( .A0(n23), .A1(n27), .B0(n31), .B1(n5), .Y(out[2]) );
  AOI31X4 U10 ( .A0(n3), .A1(n4), .A2(n5), .B0(n31), .Y(n38) );
  OAI2BB2X1 U11 ( .B0(n31), .B1(n4), .A0N(n33), .A1N(n31), .Y(out[3]) );
  OAI2BB2X2 U12 ( .B0(n31), .B1(n6), .A0N(in[1]), .A1N(n31), .Y(out[1]) );
  CLKINVX4 U13 ( .A(n23), .Y(n28) );
  BUFX2 U14 ( .A(in[4]), .Y(n23) );
  AO21XL U15 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKBUFX1TH U17 ( .A(out[6]), .Y(out[4]) );
  CLKBUFX1TH U18 ( .A(out[6]), .Y(out[5]) );
  CLKBUFX1TH U19 ( .A(in[0]), .Y(out[0]) );
  NOR2BXLTH U20 ( .AN(n6), .B(in[0]), .Y(n3) );
  NAND2XLTH U21 ( .A(n8), .B(n27), .Y(n7) );
  CLKINVX40 U16 ( .A(n28), .Y(n30) );
  CLKINVX40 U22 ( .A(n30), .Y(n31) );
  CLKBUFX40 U23 ( .A(n34), .Y(n32) );
  CLKBUFX40 U24 ( .A(in[3]), .Y(n33) );
  DLY1X1TH U25 ( .A(n37), .Y(n34) );
  CLKINVX40 U26 ( .A(n38), .Y(n35) );
  CLKINVX40 U27 ( .A(n35), .Y(out[6]) );
  XOR2X1 U28 ( .A(n7), .B(n33), .Y(n37) );
  CLKINVX40 U29 ( .A(n32), .Y(n4) );
endmodule


module sm_tc_28 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  AOI31X2TH U2 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2X3TH U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVXLTH U4 ( .A(out[4]), .Y(n18) );
  OAI2BB2X1TH U5 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  OAI2BB2X1TH U6 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U7 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U8 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U9 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U10 ( .A(n8), .B(n21), .Y(n7) );
  CLKINVX2TH U11 ( .A(in[4]), .Y(n22) );
  CLKINVX1TH U12 ( .A(n18), .Y(out[5]) );
  CLKINVX1TH U13 ( .A(in[2]), .Y(n21) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI22X1TH U15 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  XNOR2X1TH U16 ( .A(n21), .B(n8), .Y(n5) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_7_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR3X2 U3 ( .A(A[6]), .B(n3), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
  CLKINVX40 U5 ( .A(B[6]), .Y(n3) );
endmodule


module add_7_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n4, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, n1, n2;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry_6_), .Y(n4) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2])
         );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4])
         );
  ADDFX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry_2_), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKINVX40 U3 ( .A(n4), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_7_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_7_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
endmodule


module add_7_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, n1;

  ADDFHXLTH U1_5 ( .A(B[5]), .B(A[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(B[4]), .B(A[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  ADDFHX2TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  ADDFHXLTH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry_2_), .S(SUM[1]) );
  XOR3XL U1_6 ( .A(A[6]), .B(B[6]), .C(carry_6_), .Y(SUM[6]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_7_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_7 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;

  add_7_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n25, n26, n21, 
        temp1_0_}), .B({n24, in2[5:0]}), .SUM(out3) );
  add_7_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, n27, temp2_0_}), .B(in), .SUM(out1) );
  add_7_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n25, n26, n21, 
        temp1_0_}), .B({in3[6:5], n22, n28, n19, n20, in3[0]}), .SUM(out2) );
  add_7_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n25, n26, n21, 
        temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, n27, 
        temp2_0_}), .SUM(out) );
  add_7_DW01_add_4 add_30 ( .A({n23, in2[5:0]}), .B({in3[6:5], n22, n28, n19, 
        n20, in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_7_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2 U1 ( .A(in3[2]), .Y(n19) );
  CLKBUFX40 U2 ( .A(in3[1]), .Y(n20) );
  CLKBUFX40 U3 ( .A(temp1_1_), .Y(n21) );
  CLKBUFX40 U4 ( .A(in3[4]), .Y(n22) );
  DLY1X1TH U5 ( .A(in2[6]), .Y(n23) );
  DLY1X1TH U6 ( .A(in2[6]), .Y(n24) );
  CLKBUFX40 U13 ( .A(temp1_3_), .Y(n25) );
  CLKBUFX40 U14 ( .A(temp1_2_), .Y(n26) );
  CLKBUFX40 U15 ( .A(temp2_1_), .Y(n27) );
  CLKBUFX40 U16 ( .A(in3[3]), .Y(n28) );
endmodule


module tc_sm_31 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n25, n26, n28, n29, n30, n31, n32,
         n34, n35;

  BUFX3 U3 ( .A(in[6]), .Y(n25) );
  INVXLTH U4 ( .A(in[6]), .Y(n26) );
  NOR3X1TH U5 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U6 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U7 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U8 ( .A(in[2]), .Y(n31) );
  XNOR2XLTH U9 ( .A(n31), .B(n11), .Y(n10) );
  NOR2XLTH U10 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U11 ( .A0(in[4]), .A1(n35), .A2(in[5]), .B0(n13), .B1(n28), .B2(
        n29), .Y(n8) );
  INVXLTH U12 ( .A(in[5]), .Y(n28) );
  INVXLTH U13 ( .A(in[4]), .Y(n29) );
  CLKINVX1TH U14 ( .A(in[3]), .Y(n30) );
  CLKBUFX1TH U15 ( .A(n35), .Y(out[4]) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n12), .B0(n35), .B1(n32), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U18 ( .A0(n26), .A1(n10), .B0(n35), .B1(n31), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U19 ( .A0(n9), .A1(n30), .B0(n35), .Y(n7) );
  OAI211XLTH U20 ( .A0(n35), .A1(n30), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U21 ( .A0N(n30), .A1N(n9), .B0(n35), .Y(n13) );
  CLKINVX40 U22 ( .A(n25), .Y(n34) );
  CLKINVX40 U23 ( .A(n34), .Y(n35) );
endmodule


module tc_sm_30 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17, n18;

  INVXLTH U3 ( .A(in[6]), .Y(n15) );
  OAI221XLTH U4 ( .A0(n15), .A1(n8), .B0(in[6]), .B1(n17), .C0(n6), .Y(out[2])
         );
  OAI211XLTH U5 ( .A0(in[6]), .A1(n16), .B0(n5), .C0(n6), .Y(out[3]) );
  NOR3X1TH U6 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  OAI221XLTH U7 ( .A0(n15), .A1(n10), .B0(in[6]), .B1(n18), .C0(n6), .Y(out[1]) );
  OAI21BX1TH U8 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n12) );
  NAND2XL U9 ( .A(in[6]), .B(n11), .Y(n13) );
  OAI2B11X2TH U10 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  AND2X8 U11 ( .A(n13), .B(n12), .Y(n6) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  XOR2XLTH U13 ( .A(in[0]), .B(n18), .Y(n10) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  OAI21XLTH U15 ( .A0(n7), .A1(n16), .B0(in[6]), .Y(n5) );
  INVXLTH U16 ( .A(in[3]), .Y(n16) );
  INVXLTH U17 ( .A(in[1]), .Y(n18) );
  INVXLTH U18 ( .A(in[2]), .Y(n17) );
  XOR2XLTH U19 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n9) );
endmodule


module tc_sm_29 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n21, n23, n24, n25, n26, n28;

  OAI2B11X1TH U4 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OAI211XLTH U5 ( .A0(in[6]), .A1(n24), .B0(n5), .C0(n6), .Y(out[3]) );
  INVXLTH U6 ( .A(in[6]), .Y(n23) );
  AOI2BB1X1TH U7 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  OAI221XLTH U8 ( .A0(n23), .A1(n8), .B0(in[6]), .B1(n25), .C0(n6), .Y(out[2])
         );
  OAI221XLTH U9 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n26), .C0(n6), .Y(out[1]) );
  NAND2BXLTH U10 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  CLKAND2X2 U11 ( .A(in[6]), .B(n11), .Y(n21) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U14 ( .A(in[2]), .Y(n25) );
  XOR2XLTH U15 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n9) );
  XOR2XLTH U17 ( .A(in[0]), .B(n26), .Y(n10) );
  INVXLTH U18 ( .A(in[1]), .Y(n26) );
  OAI21XLTH U19 ( .A0(n7), .A1(n24), .B0(in[6]), .Y(n5) );
  INVXLTH U20 ( .A(in[3]), .Y(n24) );
  OR2X8 U3 ( .A(n21), .B(n12), .Y(n28) );
  CLKINVX40 U21 ( .A(n28), .Y(n6) );
endmodule


module tc_sm_28 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n20, n21, n22, n23, n24, n25;

  BUFX10 U3 ( .A(n8), .Y(n18) );
  OAI211XL U4 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n18), .Y(out[3]) );
  OAI221X2 U5 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n18), .Y(out[2])
         );
  OAI221XL U6 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n18), .Y(out[1])
         );
  OAI2BB1X4 U7 ( .A0N(n23), .A1N(n9), .B0(in[6]), .Y(n13) );
  INVXLTH U8 ( .A(in[6]), .Y(n20) );
  CLKINVX1TH U9 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U11 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U13 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U15 ( .A(in[2]), .Y(n24) );
  OAI21XLTH U16 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  INVX2 U19 ( .A(in[5]), .Y(n21) );
  OAI33X4 U20 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n21), .B2(
        n22), .Y(n8) );
  INVXL U21 ( .A(in[4]), .Y(n22) );
endmodule


module total_3_test_40 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n63, w5_4_, n9, n10, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_31 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_30 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_29 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_28 sm_tc_4 ( .out(in1), .in(in) );
  add_7 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), .in2(
        b1), .in3(c1), .in(in1) );
  tc_sm_31 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_30 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_29 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_28 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n59), .CK(clk), .RN(n9), 
        .Q(up3[4]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n54), .CK(clk), .RN(n10), 
        .Q(h) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n58), .CK(clk), .RN(n9), 
        .Q(up3[3]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n59), .CK(clk), .RN(n9), 
        .Q(up3[2]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n50), .CK(clk), .RN(n9), 
        .Q(up2[0]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n50), .CK(clk), .RN(n9), 
        .Q(up3[0]) );
  SDFFRQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n53), .CK(clk), .RN(n9), 
        .Q(up1[4]) );
  SDFFRQX2TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n58), .CK(clk), .RN(n9), .Q(
        up1[0]) );
  SDFFRQX1TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n49), .CK(clk), .RN(n10), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n56), .CK(clk), .RN(n9), 
        .Q(n63) );
  SDFFRQX1 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n49), .CK(clk), .RN(n9), 
        .Q(up2[1]) );
  SDFFRQX1 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n56), .CK(clk), .RN(n9), 
        .Q(up2[2]) );
  SDFFRQX1 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n54), .CK(clk), .RN(n9), 
        .Q(up2[3]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n10) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n9) );
  SDFFRHQX8 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n57), .CK(clk), .RN(n9), 
        .Q(up1[1]) );
  SDFFRHQX8 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n53), .CK(clk), .RN(n9), 
        .Q(up1[2]) );
  SDFFRHQX8 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n57), .CK(clk), .RN(n10), 
        .Q(up1[3]) );
  DLY1X1TH U37 ( .A(n63), .Y(up3[1]) );
  INVXLTH U38 ( .A(n51), .Y(n49) );
  INVXLTH U39 ( .A(n52), .Y(n50) );
  DLY1X1TH U40 ( .A(n55), .Y(n51) );
  DLY1X1TH U41 ( .A(n55), .Y(n52) );
  INVXLTH U42 ( .A(n52), .Y(n53) );
  INVXLTH U43 ( .A(n51), .Y(n54) );
  INVXLTH U44 ( .A(test_se), .Y(n55) );
  INVXLTH U45 ( .A(n52), .Y(n56) );
  INVXLTH U46 ( .A(n51), .Y(n57) );
  INVXLTH U47 ( .A(n52), .Y(n58) );
  INVXLTH U48 ( .A(n51), .Y(n59) );
endmodule


module sm_tc_27 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n21, n25, n26;

  OAI2BB2X1 U2 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  AOI31X2 U3 ( .A0(n3), .A1(n4), .A2(n5), .B0(n26), .Y(out[4]) );
  OAI2BB2X1 U4 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n26), .Y(out[1]) );
  INVX6 U6 ( .A(n21), .Y(n26) );
  BUFX6 U7 ( .A(in[4]), .Y(n21) );
  NOR2X2 U8 ( .A(in[1]), .B(in[0]), .Y(n8) );
  XNOR2X1TH U9 ( .A(n25), .B(n8), .Y(n5) );
  BUFX2TH U10 ( .A(in[0]), .Y(out[0]) );
  INVX2TH U11 ( .A(in[2]), .Y(n25) );
  CLKNAND2X2TH U12 ( .A(n8), .B(n25), .Y(n7) );
  AO21X4 U13 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  XNOR2X2TH U14 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[6]) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  AO2B2BX4 U5 ( .A0(n26), .A1N(n25), .B0(n21), .B1N(n5), .Y(out[2]) );
endmodule


module sm_tc_26 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n25, n26, n27, n28, n29;

  AOI31X2TH U3 ( .A0(n6), .A1(n27), .A2(n3), .B0(n25), .Y(out[4]) );
  INVX2TH U4 ( .A(in[4]), .Y(n25) );
  CLKBUFX1TH U5 ( .A(in[0]), .Y(out[0]) );
  XNOR2X2TH U6 ( .A(n26), .B(n8), .Y(n4) );
  OAI22X1TH U7 ( .A0(in[4]), .A1(n26), .B0(n25), .B1(n4), .Y(out[2]) );
  INVX2TH U8 ( .A(in[2]), .Y(n26) );
  XNOR2X2TH U10 ( .A(n7), .B(in[3]), .Y(n3) );
  NOR2BXLTH U12 ( .AN(n5), .B(in[0]), .Y(n6) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[6]) );
  NAND2XLTH U15 ( .A(n8), .B(n26), .Y(n7) );
  AO21XLTH U16 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n5) );
  XNOR2X2TH U2 ( .A(n26), .B(n8), .Y(n27) );
  AO2B2X4 U9 ( .B0(in[1]), .B1(n25), .A0(n29), .A1N(n5), .Y(out[1]) );
  OR2X8 U11 ( .A(in[1]), .B(in[0]), .Y(n28) );
  CLKINVX40 U17 ( .A(n28), .Y(n8) );
  AO2B2BX4 U18 ( .A0(n29), .A1N(n3), .B0(in[3]), .B1N(n29), .Y(out[3]) );
  CLKINVX40 U19 ( .A(n25), .Y(n29) );
endmodule


module sm_tc_25 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n29, n30, n33, n34, n35;

  OAI2BB2X2 U5 ( .B0(n30), .B1(n6), .A0N(in[1]), .A1N(n30), .Y(out[1]) );
  OAI22XL U3 ( .A0(in[4]), .A1(n33), .B0(n30), .B1(n5), .Y(out[2]) );
  CLKINVX1TH U6 ( .A(in[2]), .Y(n29) );
  NAND2X1TH U7 ( .A(n8), .B(n33), .Y(n7) );
  INVX2TH U8 ( .A(in[4]), .Y(n30) );
  OAI2BB2X1TH U9 ( .B0(n30), .B1(n4), .A0N(in[3]), .A1N(n30), .Y(out[3]) );
  AO21X1TH U10 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  XNOR2X2TH U11 ( .A(n7), .B(in[3]), .Y(n4) );
  AOI31X2TH U12 ( .A0(n3), .A1(n4), .A2(n34), .B0(n30), .Y(out[4]) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[6]) );
  BUFX2TH U16 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX40 U2 ( .A(n29), .Y(n33) );
  XOR2X1 U4 ( .A(n33), .B(n35), .Y(n34) );
  OR2X8 U17 ( .A(in[1]), .B(in[0]), .Y(n35) );
  CLKINVX40 U18 ( .A(n35), .Y(n8) );
  XOR2X1 U19 ( .A(n33), .B(n35), .Y(n5) );
endmodule


module sm_tc_24 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  OAI22X1TH U2 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  XNOR2X1TH U3 ( .A(n7), .B(in[3]), .Y(n4) );
  INVXLTH U4 ( .A(n18), .Y(out[6]) );
  NOR2X3TH U5 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVXLTH U6 ( .A(n18), .Y(out[5]) );
  OAI2BB2X1TH U7 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  AO21X1TH U8 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  XNOR2X1TH U9 ( .A(n21), .B(n8), .Y(n5) );
  CLKINVX1TH U10 ( .A(in[2]), .Y(n21) );
  NAND2XLTH U11 ( .A(n8), .B(n21), .Y(n7) );
  CLKINVX2TH U12 ( .A(in[4]), .Y(n22) );
  INVXLTH U13 ( .A(out[4]), .Y(n18) );
  AOI31X4TH U14 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2BB2X1TH U16 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  CLKBUFX1TH U17 ( .A(in[0]), .Y(out[0]) );
endmodule


module add_6_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_6_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8;
  wire   [6:2] carry;

  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n5), .CO(carry[2]), .S(SUM[1]) );
  ADDFX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  NAND2XL U1 ( .A(carry[4]), .B(n7), .Y(n2) );
  NAND2X1TH U2 ( .A(n7), .B(B[4]), .Y(n4) );
  CLKXOR2X1TH U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND3X2 U6 ( .A(n2), .B(n3), .C(n4), .Y(carry[5]) );
  AND2XLTH U7 ( .A(B[0]), .B(A[0]), .Y(n5) );
  XNOR2X1 U3 ( .A(n6), .B(carry[4]), .Y(SUM[4]) );
  XNOR2X4 U5 ( .A(B[4]), .B(n7), .Y(n6) );
  CLKBUFX40 U8 ( .A(A[4]), .Y(n7) );
  AND2X8 U9 ( .A(carry[4]), .B(B[4]), .Y(n8) );
  CLKINVX40 U10 ( .A(n8), .Y(n3) );
endmodule


module add_6_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_6_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n14, n2, n4, n7, n8, n9, n10, n11, n12;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n4), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKAND2X2TH U1 ( .A(n7), .B(n8), .Y(n9) );
  XNOR2X4 U2 ( .A(n9), .B(carry[6]), .Y(n14) );
  AND2XLTH U3 ( .A(B[0]), .B(A[0]), .Y(n4) );
  INVXLTH U4 ( .A(A[6]), .Y(n11) );
  CLKINVX1TH U5 ( .A(n2), .Y(SUM[0]) );
  XNOR2XLTH U6 ( .A(B[0]), .B(A[0]), .Y(n2) );
  NAND2XLTH U7 ( .A(n10), .B(A[6]), .Y(n8) );
  NAND2XLTH U8 ( .A(B[6]), .B(n11), .Y(n7) );
  INVXLTH U9 ( .A(B[6]), .Y(n10) );
  CLKINVX40 U10 ( .A(n14), .Y(n12) );
  CLKINVX40 U11 ( .A(n12), .Y(SUM[6]) );
endmodule


module add_6_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n6, n1, n2, n3, n4;
  wire   [6:2] carry;

  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(n6) );
  ADDFHX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR3X4 U3 ( .A(carry[3]), .B(B[3]), .C(A[3]), .Y(SUM[3]) );
  NAND2X8 U4 ( .A(carry[3]), .B(B[3]), .Y(n2) );
  NAND2X8 U5 ( .A(carry[3]), .B(A[3]), .Y(n3) );
  NAND2X8 U6 ( .A(B[3]), .B(A[3]), .Y(n4) );
  NAND3X8 U7 ( .A(n2), .B(n3), .C(n4), .Y(carry[4]) );
  CLKBUFX40 U8 ( .A(n6), .Y(SUM[5]) );
endmodule


module add_6_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n3, n1;
  wire   [6:2] carry;

  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(n3) );
  ADDFX1 U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X3TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  CLKBUFX40 U3 ( .A(n3), .Y(SUM[3]) );
endmodule


module add_6 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n22, n23, n24, n25, n26;

  add_6_DW01_add_0 add_34 ( .A({n25, temp1_5_, temp1_4_, temp1_3_, temp1_2_, 
        n22, temp1_0_}), .B({in2[6:3], n24, in2[1:0]}), .SUM(out3) );
  add_6_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_6_DW01_add_2 add_32 ( .A({n25, temp1_5_, temp1_4_, temp1_3_, temp1_2_, 
        n22, temp1_0_}), .B({in3[6:4], n26, n23, in3[1:0]}), .SUM(out2) );
  add_6_DW01_add_3 add_31 ( .A({n25, temp1_5_, temp1_4_, temp1_3_, temp1_2_, 
        n22, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_6_DW01_add_4 add_30 ( .A({in2[6:3], n24, in2[1:0]}), .B({in3[6:4], n26, 
        n23, in3[1:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}) );
  add_6_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2 U1 ( .A(temp1_1_), .Y(n22) );
  BUFX2TH U2 ( .A(in3[2]), .Y(n23) );
  CLKBUFX40 U3 ( .A(in2[2]), .Y(n24) );
  CLKBUFX40 U4 ( .A(temp1_6_), .Y(n25) );
  CLKBUFX40 U5 ( .A(in3[3]), .Y(n26) );
endmodule


module tc_sm_27 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n28) );
  XNOR2XLTH U7 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(in[6]), .Y(n24) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXLTH U11 ( .A(in[5]), .Y(n25) );
  INVXLTH U12 ( .A(in[4]), .Y(n26) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n27) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI21XLTH U16 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  OAI221XLTH U17 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U18 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(
        out[2]) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_26 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n36, n37, n38, n39, n41, n42;

  NAND2BX2 U4 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  INVXLTH U5 ( .A(in[6]), .Y(n36) );
  OAI221X2TH U7 ( .A0(n36), .A1(n8), .B0(in[6]), .B1(n38), .C0(n6), .Y(out[2])
         );
  OAI2B11X4 U9 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OAI221X2TH U10 ( .A0(n36), .A1(n10), .B0(in[6]), .B1(n39), .C0(n6), .Y(
        out[1]) );
  OAI211X2TH U11 ( .A0(in[6]), .A1(n37), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI21XLTH U12 ( .A0(n7), .A1(n37), .B0(in[6]), .Y(n5) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  INVXLTH U14 ( .A(in[2]), .Y(n38) );
  XOR2XLTH U15 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n9) );
  INVXLTH U17 ( .A(in[3]), .Y(n37) );
  CLKBUFX1TH U18 ( .A(in[6]), .Y(out[4]) );
  XOR2XLTH U19 ( .A(in[0]), .B(n39), .Y(n10) );
  INVXLTH U20 ( .A(in[1]), .Y(n39) );
  NOR2X8 U3 ( .A(n41), .B(n42), .Y(n6) );
  CLKAND2X12 U6 ( .A(in[6]), .B(n11), .Y(n41) );
  AOI2BB1X4 U8 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n42) );
endmodule


module tc_sm_25 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n18, n19, n20, n21, n22, n24, n25, n26,
         n27, n28, n29;

  CLKINVX4TH U3 ( .A(n18), .Y(n8) );
  AOI33X4 U4 ( .A0(n26), .A1(n19), .A2(n25), .B0(n20), .B1(in[5]), .B2(in[4]), 
        .Y(n18) );
  CLKINVX40 U5 ( .A(in[6]), .Y(n19) );
  AOI21BX2 U6 ( .A0(n27), .A1(n9), .B0N(in[6]), .Y(n20) );
  INVX2TH U7 ( .A(in[5]), .Y(n25) );
  OAI221XLTH U8 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n8), .Y(out[1]) );
  OAI211XLTH U9 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OR3XLTH U10 ( .A(n21), .B(n22), .C(n18), .Y(out[2]) );
  NAND2BXLTH U11 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  NOR2XLTH U12 ( .A(n24), .B(n10), .Y(n21) );
  NOR2XLTH U13 ( .A(in[6]), .B(n28), .Y(n22) );
  INVXLTH U14 ( .A(in[6]), .Y(n24) );
  CLKINVX1TH U15 ( .A(in[3]), .Y(n27) );
  NOR3X1TH U16 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U17 ( .A(in[4]), .Y(n26) );
  INVXLTH U18 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U20 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U22 ( .A(in[2]), .Y(n28) );
  CLKBUFX1TH U23 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U24 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
endmodule


module tc_sm_24 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n23, n24, n25, n27, n28, n29,
         n30, n31, n32;

  OAI211XL U3 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221XL U5 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[2])
         );
  OAI221XL U7 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[1])
         );
  INVXLTH U8 ( .A(in[6]), .Y(n20) );
  INVX2TH U9 ( .A(in[5]), .Y(n21) );
  CLKINVX1TH U11 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U12 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U14 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[2]), .Y(n24) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  CLKBUFX1TH U18 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U19 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI21XLTH U21 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  DLY1X1TH U4 ( .A(in[4]), .Y(n27) );
  AOI33X4 U6 ( .A0(n29), .A1(n30), .A2(n21), .B0(n32), .B1(n31), .B2(in[4]), 
        .Y(n28) );
  CLKINVX40 U10 ( .A(n28), .Y(n8) );
  CLKINVX40 U13 ( .A(n27), .Y(n29) );
  CLKINVX40 U22 ( .A(in[6]), .Y(n30) );
  CLKINVX40 U23 ( .A(n21), .Y(n31) );
  AOI21BX4 U24 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n32) );
endmodule


module total_3_test_41 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n6, n7, n8, n43, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_27 sm_tc_1 ( .out(a1), .in({a[4], n43, a[2:0]}) );
  sm_tc_26 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_25 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_24 sm_tc_4 ( .out(in1), .in(in) );
  add_6 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1({a1[6:1], 
        n6}), .in2(b1), .in3(c1), .in(in1) );
  tc_sm_27 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_26 tc_sm_2 ( .out(w6), .in({n59, w66[5:0]}) );
  tc_sm_25 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_24 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n58), .CK(clk), .RN(n7), 
        .Q(up3[3]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n49), .CK(clk), .RN(n7), 
        .Q(up2[3]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n57), .CK(clk), .RN(n7), 
        .Q(up3[4]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n55), .CK(clk), .RN(n7), .Q(
        up1[0]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n56), .CK(clk), .RN(n8), 
        .Q(up1[3]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n53), .CK(clk), .RN(n8), .Q(
        h) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n52), .CK(clk), .RN(n7), 
        .Q(up3[2]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n53), .CK(clk), .RN(n7), 
        .Q(up2[0]) );
  SDFFRQXLTH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n48), .CK(clk), .RN(n8), 
        .Q(up1[1]) );
  SDFFRQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n49), .CK(clk), .RN(n7), 
        .Q(up1[4]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n52), .CK(clk), .RN(n7), 
        .Q(up2[4]) );
  SDFFRQX1TH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n56), .CK(clk), .RN(n7), 
        .Q(up3[0]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n58), .CK(clk), .RN(n7), 
        .Q(up2[2]) );
  CLKBUFX2TH U3 ( .A(a1[0]), .Y(n6) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n7) );
  CLKBUFX1TH U5 ( .A(rst), .Y(n8) );
  SDFFRX4 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n57), .CK(clk), .RN(n7), 
        .Q(up1[2]) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n55), .CK(clk), .RN(n7), 
        .Q(up2[1]) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n48), .CK(clk), .RN(n7), 
        .Q(up3[1]) );
  CLKBUFX40 U38 ( .A(a[3]), .Y(n43) );
  INVXLTH U39 ( .A(n50), .Y(n48) );
  INVXLTH U40 ( .A(n51), .Y(n49) );
  DLY1X1TH U41 ( .A(n54), .Y(n50) );
  DLY1X1TH U42 ( .A(n54), .Y(n51) );
  INVXLTH U43 ( .A(n51), .Y(n52) );
  INVXLTH U44 ( .A(n50), .Y(n53) );
  INVXLTH U45 ( .A(test_se), .Y(n54) );
  INVXLTH U46 ( .A(n51), .Y(n55) );
  INVXLTH U47 ( .A(n50), .Y(n56) );
  INVXLTH U48 ( .A(n51), .Y(n57) );
  INVXLTH U49 ( .A(n50), .Y(n58) );
  CLKBUFX40 U50 ( .A(w66[6]), .Y(n59) );
endmodule


module sm_tc_23 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n24, n25, n28, n29, n30;

  XNOR2X2 U3 ( .A(n24), .B(n8), .Y(n5) );
  OAI22XL U4 ( .A0(in[4]), .A1(n24), .B0(n25), .B1(n5), .Y(out[2]) );
  INVX2TH U6 ( .A(in[2]), .Y(n24) );
  CLKBUFX2 U7 ( .A(in[0]), .Y(out[0]) );
  AO21X4 U8 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2XLTH U9 ( .B0(n25), .B1(n4), .A0N(in[3]), .A1N(n25), .Y(out[3]) );
  INVX4TH U11 ( .A(in[4]), .Y(n25) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[6]) );
  AOI31X2TH U13 ( .A0(n3), .A1(n4), .A2(n5), .B0(n25), .Y(out[4]) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2X4 U16 ( .B0(n25), .B1(n6), .A0N(in[1]), .A1N(n25), .Y(out[1]) );
  NAND2BX8 U2 ( .AN(in[1]), .B(n29), .Y(n28) );
  CLKINVX40 U5 ( .A(n28), .Y(n8) );
  CLKINVX40 U10 ( .A(in[0]), .Y(n29) );
  XOR2X1 U17 ( .A(n30), .B(in[3]), .Y(n4) );
  CLKAND2X12 U18 ( .A(n8), .B(n24), .Y(n30) );
endmodule


module sm_tc_22 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n21, n22, n25;

  OAI2BB2X4 U2 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  NOR2X4 U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  BUFX6 U4 ( .A(in[4]), .Y(n17) );
  AO21X1 U7 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  AOI31X2TH U9 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  CLKBUFX1TH U10 ( .A(out[4]), .Y(out[5]) );
  CLKINVX1TH U11 ( .A(in[2]), .Y(n21) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[6]) );
  CLKNAND2X4 U13 ( .A(n8), .B(n21), .Y(n7) );
  XNOR2X2TH U14 ( .A(n7), .B(in[3]), .Y(n4) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  BUFX2TH U16 ( .A(in[0]), .Y(out[0]) );
  INVX3 U17 ( .A(n17), .Y(n22) );
  OAI2B2X2 U5 ( .A1N(in[3]), .A0(n17), .B0(n22), .B1(n4), .Y(out[3]) );
  OAI2B2X2 U6 ( .A1N(n17), .A0(n5), .B0(n17), .B1(n21), .Y(out[2]) );
  XOR2X1 U8 ( .A(n21), .B(n25), .Y(n5) );
  CLKINVX40 U18 ( .A(n8), .Y(n25) );
endmodule


module sm_tc_21 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n28, n29, n32, n33, n34, n35;

  INVX2 U2 ( .A(in[4]), .Y(n29) );
  OAI2BB2XL U3 ( .B0(n35), .B1(n4), .A0N(in[3]), .A1N(n35), .Y(out[3]) );
  AO21X2 U5 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI22X2 U6 ( .A0(n34), .A1(n28), .B0(n35), .B1(n5), .Y(out[2]) );
  AOI31X2 U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n35), .Y(out[4]) );
  CLKBUFX1TH U8 ( .A(out[4]), .Y(out[6]) );
  INVX1TH U9 ( .A(in[2]), .Y(n28) );
  XNOR2X2TH U10 ( .A(n7), .B(in[3]), .Y(n4) );
  XNOR2X1TH U12 ( .A(n28), .B(n8), .Y(n5) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  BUFX2TH U15 ( .A(in[0]), .Y(out[0]) );
  NAND2XLTH U16 ( .A(n8), .B(n28), .Y(n7) );
  OR2X8 U4 ( .A(in[1]), .B(in[0]), .Y(n32) );
  CLKINVX40 U11 ( .A(n32), .Y(n8) );
  AO2B2X4 U17 ( .B0(in[1]), .B1(n35), .A0(n34), .A1N(n6), .Y(out[1]) );
  CLKBUFX40 U18 ( .A(n29), .Y(n33) );
  CLKINVX40 U19 ( .A(n33), .Y(n34) );
  CLKINVX40 U20 ( .A(n34), .Y(n35) );
endmodule


module sm_tc_20 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  AO21X1TH U2 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X3TH U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI2BB2X1TH U4 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U5 ( .A(in[0]), .Y(out[0]) );
  CLKINVX1TH U6 ( .A(in[2]), .Y(n21) );
  CLKINVX2TH U7 ( .A(in[4]), .Y(n22) );
  AOI31X2TH U8 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U9 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U10 ( .A(out[4]), .Y(n18) );
  INVXLTH U11 ( .A(n18), .Y(out[5]) );
  OAI22X1TH U12 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  OAI2BB2X1TH U13 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  INVXLTH U14 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U15 ( .A(n21), .B(n8), .Y(n5) );
  XNOR2X1TH U16 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U17 ( .A(n8), .B(n21), .Y(n7) );
endmodule


module add_5_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKAND2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_5_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n4, n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n4) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  CLKINVX40 U3 ( .A(n4), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_5_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X4TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_5_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n3, n4;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n3) );
  CLKINVX1TH U2 ( .A(n1), .Y(SUM[0]) );
  XNOR2XLTH U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U4 ( .A(n4), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKINVX40 U5 ( .A(A[6]), .Y(n4) );
endmodule


module add_5_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [6:2] carry;

  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX4 U1_2 ( .A(carry[2]), .B(B[2]), .CI(A[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKXOR2X2 U1 ( .A(A[5]), .B(B[5]), .Y(n6) );
  NAND3X2 U2 ( .A(n3), .B(n4), .C(n5), .Y(carry[4]) );
  NAND2XLTH U3 ( .A(B[3]), .B(A[3]), .Y(n3) );
  NAND2XLTH U4 ( .A(A[3]), .B(carry[3]), .Y(n5) );
  XOR2X3 U5 ( .A(n2), .B(B[3]), .Y(SUM[3]) );
  CLKXOR2X2TH U6 ( .A(n6), .B(carry[5]), .Y(SUM[5]) );
  CLKNAND2X2TH U7 ( .A(carry[5]), .B(B[5]), .Y(n7) );
  NAND2XL U8 ( .A(carry[5]), .B(A[5]), .Y(n8) );
  XOR2X1TH U9 ( .A(carry[3]), .B(A[3]), .Y(n2) );
  NAND2XLTH U10 ( .A(B[5]), .B(A[5]), .Y(n9) );
  NAND3X2TH U11 ( .A(n7), .B(n8), .C(n9), .Y(carry[6]) );
  NAND2XLTH U12 ( .A(B[3]), .B(carry[3]), .Y(n4) );
  CLKXOR2X2TH U13 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U14 ( .A(A[0]), .B(B[0]), .Y(n1) );
endmodule


module add_5_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2TH U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_5 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n20, n21, n22, n23;

  add_5_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n23, temp1_0_}), .B(in2), .SUM(out3) );
  add_5_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_5_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n23, temp1_0_}), .B({in3[6:4], n21, in3[2:0]}), .SUM(out2)
         );
  add_5_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n23, temp1_0_}), .B({temp2_6_, n22, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_5_DW01_add_4 add_30 ( .A(in2), .B({in3[6:4], n21, in3[2:0]}), .SUM({
        temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_})
         );
  add_5_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  INVX3 U1 ( .A(in3[3]), .Y(n20) );
  INVX4 U2 ( .A(n20), .Y(n21) );
  CLKBUFX1TH U3 ( .A(temp2_5_), .Y(n22) );
  CLKBUFX40 U4 ( .A(temp1_1_), .Y(n23) );
endmodule


module tc_sm_23 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29;

  CLKBUFX1 U3 ( .A(in[6]), .Y(out[4]) );
  NOR3X1TH U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U5 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U6 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U7 ( .A(in[2]), .Y(n28) );
  XNOR2XLTH U8 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXLTH U11 ( .A(in[5]), .Y(n25) );
  INVXLTH U12 ( .A(in[4]), .Y(n26) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n27) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n24) );
  OAI221XLTH U16 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_22 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n25, n26, n27, n29, n30, n31, n32;

  NAND3XL U3 ( .A(n26), .B(n27), .C(n6), .Y(out[2]) );
  OA21XL U4 ( .A0(in[6]), .A1(n30), .B0(n5), .Y(n25) );
  NAND2XLTH U5 ( .A(n25), .B(n6), .Y(out[3]) );
  OAI21X1 U6 ( .A0(n7), .A1(n30), .B0(in[6]), .Y(n5) );
  AOI21X8 U7 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n6) );
  INVXL U8 ( .A(in[6]), .Y(n29) );
  OR2X2 U9 ( .A(n29), .B(n8), .Y(n26) );
  XOR2XLTH U10 ( .A(in[2]), .B(n9), .Y(n8) );
  CLKBUFX1TH U11 ( .A(in[6]), .Y(out[4]) );
  OAI221X1TH U12 ( .A0(n29), .A1(n10), .B0(in[6]), .B1(n32), .C0(n6), .Y(
        out[1]) );
  OR2XL U13 ( .A(in[6]), .B(n31), .Y(n27) );
  OAI2B11X2 U14 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  AOI2BB1X4 U15 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  NOR3X1TH U16 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  XOR2XLTH U17 ( .A(in[0]), .B(n32), .Y(n10) );
  INVXLTH U18 ( .A(in[1]), .Y(n32) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  INVXLTH U20 ( .A(in[2]), .Y(n31) );
  NOR2XLTH U21 ( .A(in[0]), .B(in[1]), .Y(n9) );
  INVXLTH U22 ( .A(in[3]), .Y(n30) );
endmodule


module tc_sm_21 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n21, n22, n23, n24, n26;

  AOI2BB1X2TH U4 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n12) );
  OAI2B11X1TH U5 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  NOR3X1TH U6 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  INVXLTH U7 ( .A(in[2]), .Y(n23) );
  XOR2XLTH U8 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI211XLTH U10 ( .A0(in[6]), .A1(n22), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI21XLTH U11 ( .A0(n7), .A1(n22), .B0(in[6]), .Y(n5) );
  INVXLTH U12 ( .A(in[3]), .Y(n22) );
  XOR2XLTH U13 ( .A(in[0]), .B(n24), .Y(n10) );
  INVXLTH U14 ( .A(in[1]), .Y(n24) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U16 ( .A(in[6]), .Y(n21) );
  OAI221XLTH U17 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n24), .C0(n6), .Y(
        out[1]) );
  OAI221XLTH U18 ( .A0(n21), .A1(n8), .B0(in[6]), .B1(n23), .C0(n6), .Y(out[2]) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  AO21X4 U3 ( .A0(in[6]), .A1(n11), .B0(n12), .Y(n26) );
  CLKINVX40 U20 ( .A(n26), .Y(n6) );
endmodule


module tc_sm_20 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n26, n27,
         n28;

  OAI221XL U3 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1])
         );
  OAI221XL U4 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2])
         );
  NAND2BXLTH U5 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211XLTH U6 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  CLKINVX1TH U7 ( .A(in[3]), .Y(n22) );
  INVXLTH U8 ( .A(in[4]), .Y(n21) );
  INVXLTH U9 ( .A(in[5]), .Y(n20) );
  NOR3X1TH U10 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U11 ( .A(in[6]), .Y(n19) );
  INVXLTH U12 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U14 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[2]), .Y(n23) );
  OAI21XLTH U17 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U18 ( .A(in[6]), .Y(out[4]) );
  AOI33X4 U19 ( .A0(n21), .A1(n27), .A2(n20), .B0(n28), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U20 ( .A(n26), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n27) );
  AOI21BX4 U22 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n28) );
endmodule


module total_3_test_42 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n4, n5, n44, n45, n46, n47, n48, n49, n50, n51;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_23 sm_tc_1 ( .out(a1), .in({n4, a[3:0]}) );
  sm_tc_22 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_21 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_20 sm_tc_4 ( .out(in1), .in(in) );
  add_5 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), .in2(
        b1), .in3(c1), .in(in1) );
  tc_sm_23 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_22 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_21 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_20 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n49), .CK(clk), .RN(rst), 
        .Q(up3[4]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(test_se), .CK(clk), .RN(n5), 
        .Q(up1[0]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n47), .CK(clk), .RN(n5), .Q(
        h) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(test_se), .CK(clk), .RN(
        n5), .Q(up3[3]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n47), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRQX1TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  SDFFRQXL up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up1[2]) );
  SDFFRQX1 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n45), .CK(clk), .RN(n5), 
        .Q(up2[1]) );
  SDFFRQX1 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n47), .CK(clk), .RN(n5), 
        .Q(up2[2]) );
  SDFFRQX4 up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  BUFX4 U3 ( .A(a[4]), .Y(n4) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n5) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n47), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  SDFFRX4 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n45), .CK(clk), .RN(rst), 
        .Q(up1[3]) );
  SDFFRX4 up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  DLY1X1TH U37 ( .A(n48), .Y(n44) );
  INVXLTH U38 ( .A(n44), .Y(n45) );
  INVXLTH U39 ( .A(n48), .Y(n46) );
  DLY1X1TH U40 ( .A(test_se), .Y(n47) );
  INVXLTH U41 ( .A(test_se), .Y(n48) );
  INVXLTH U42 ( .A(n44), .Y(n49) );
  INVXLTH U43 ( .A(n44), .Y(n50) );
  INVXLTH U44 ( .A(n44), .Y(n51) );
endmodule


module sm_tc_19 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n21, n22;

  OAI22X4 U2 ( .A0(n17), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  OAI2BB2X2 U3 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  AOI31X2TH U4 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  INVX18 U5 ( .A(n17), .Y(n22) );
  BUFX10 U6 ( .A(in[4]), .Y(n17) );
  INVX2 U7 ( .A(in[2]), .Y(n21) );
  XNOR2X1 U8 ( .A(n7), .B(in[3]), .Y(n4) );
  BUFX3 U9 ( .A(in[0]), .Y(out[0]) );
  CLKBUFX1TH U10 ( .A(out[4]), .Y(out[6]) );
  OAI2BB2X4 U11 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  XNOR2X4TH U12 ( .A(n21), .B(n8), .Y(n5) );
  AO21X2TH U13 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X6 U14 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  NAND2XLTH U16 ( .A(n8), .B(n21), .Y(n7) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
endmodule


module sm_tc_18 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n29, n30, n31, n35, n36;

  CLKINVX2 U2 ( .A(n36), .Y(n29) );
  INVX4 U3 ( .A(in[4]), .Y(n36) );
  XNOR2X1TH U4 ( .A(n7), .B(in[3]), .Y(n4) );
  NAND2XLTH U5 ( .A(n8), .B(n35), .Y(n7) );
  CLKBUFX1TH U6 ( .A(out[4]), .Y(out[6]) );
  AOI31X4TH U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n36), .Y(out[4]) );
  OAI2BB2X1TH U8 ( .B0(n36), .B1(n6), .A0N(in[1]), .A1N(n36), .Y(out[1]) );
  AO21X1TH U9 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X4 U10 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX2 U11 ( .A(in[2]), .Y(n35) );
  XNOR2X4TH U12 ( .A(n35), .B(n8), .Y(n5) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  OR2XLTH U15 ( .A(n29), .B(n35), .Y(n30) );
  OR2XLTH U16 ( .A(n36), .B(n5), .Y(n31) );
  NAND2X1TH U17 ( .A(n30), .B(n31), .Y(out[2]) );
  OAI2BB2X1TH U18 ( .B0(n36), .B1(n4), .A0N(in[3]), .A1N(n36), .Y(out[3]) );
  CLKBUFX1TH U19 ( .A(in[0]), .Y(out[0]) );
endmodule


module sm_tc_17 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n23, n27, n28, n31, n32;

  NOR2X4 U2 ( .A(n31), .B(out[0]), .Y(n8) );
  CLKBUFX4 U3 ( .A(in[0]), .Y(out[0]) );
  AO21XL U5 ( .A0(out[0]), .A1(n31), .B0(n8), .Y(n6) );
  XNOR2X4 U6 ( .A(n28), .B(n8), .Y(n5) );
  BUFX3 U7 ( .A(in[4]), .Y(n23) );
  OAI2BB2X4 U9 ( .B0(n27), .B1(n6), .A0N(n31), .A1N(n27), .Y(out[1]) );
  OAI22XLTH U10 ( .A0(n23), .A1(n28), .B0(n27), .B1(n5), .Y(out[2]) );
  INVX2 U11 ( .A(n23), .Y(n27) );
  AOI31X2 U12 ( .A0(n3), .A1(n4), .A2(n5), .B0(n27), .Y(out[4]) );
  CLKINVX1TH U13 ( .A(in[2]), .Y(n28) );
  NOR2BXLTH U15 ( .AN(n6), .B(out[0]), .Y(n3) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[6]) );
  AO2B2X4 U4 ( .B0(in[3]), .B1(n27), .A0(n23), .A1N(n4), .Y(out[3]) );
  CLKBUFX40 U8 ( .A(in[1]), .Y(n31) );
  XOR2X1 U14 ( .A(n32), .B(in[3]), .Y(n4) );
  CLKAND2X12 U18 ( .A(n8), .B(n28), .Y(n32) );
endmodule


module sm_tc_16 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  CLKBUFX2TH U2 ( .A(in[0]), .Y(out[0]) );
  NOR2X3 U3 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX1TH U4 ( .A(in[2]), .Y(n21) );
  AOI31X2TH U5 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U6 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U7 ( .A(n18), .Y(out[5]) );
  OAI2BB2X1TH U8 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  NAND2XLTH U9 ( .A(n8), .B(n21), .Y(n7) );
  INVXLTH U10 ( .A(n18), .Y(out[6]) );
  XNOR2X1TH U11 ( .A(n21), .B(n8), .Y(n5) );
  CLKINVX2TH U12 ( .A(in[4]), .Y(n22) );
  INVXLTH U13 ( .A(out[4]), .Y(n18) );
  OAI22X1TH U14 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  OAI2BB2X1TH U15 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  XNOR2X1TH U16 ( .A(n7), .B(in[3]), .Y(n4) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_4_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [6:2] carry;

  NAND3X2 U5 ( .A(n2), .B(n3), .C(n4), .Y(carry[5]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n5), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X2 U2 ( .A(B[0]), .B(A[0]), .Y(n5) );
  CLKNAND2X2TH U3 ( .A(n8), .B(n9), .Y(SUM[4]) );
  CLKINVX4TH U4 ( .A(n1), .Y(n6) );
  NAND2XLTH U7 ( .A(A[4]), .B(B[4]), .Y(n3) );
  CLKNAND2X2TH U8 ( .A(A[4]), .B(carry[4]), .Y(n2) );
  NAND2XLTH U9 ( .A(n6), .B(A[4]), .Y(n9) );
  NAND2XLTH U10 ( .A(n1), .B(n7), .Y(n8) );
  INVXLTH U11 ( .A(A[4]), .Y(n7) );
  CLKXOR2X2TH U12 ( .A(B[4]), .B(carry[4]), .Y(n1) );
  XNOR3X2 U6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n10) );
  CLKINVX40 U13 ( .A(n10), .Y(SUM[6]) );
  AND2X8 U14 ( .A(carry[4]), .B(B[4]), .Y(n11) );
  CLKINVX40 U15 ( .A(n11), .Y(n4) );
endmodule


module add_4_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n4, n1, n2;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n4) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  CLKINVX40 U3 ( .A(n4), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_4_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X12 U1 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  CLKXOR2X1TH U3 ( .A(B[6]), .B(A[6]), .Y(n2) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_4_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3;
  wire   [6:2] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX1 U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  DLY1X1TH U2 ( .A(n3), .Y(n2) );
  XNOR2X1 U3 ( .A(B[0]), .B(A[0]), .Y(n3) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[0]) );
endmodule


module add_4_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [6:2] carry;

  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(carry[4]), .CI(B[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  NAND2X2 U1 ( .A(n4), .B(n5), .Y(SUM[0]) );
  NAND2XLTH U2 ( .A(B[0]), .B(n3), .Y(n4) );
  NAND2XL U3 ( .A(n2), .B(A[0]), .Y(n5) );
  INVXLTH U4 ( .A(B[0]), .Y(n2) );
  INVXLTH U5 ( .A(A[0]), .Y(n3) );
  AND2XLTH U6 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_4 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         add_31_n6, add_31_n5, add_31_n4, add_31_n1, add_31_carry_2_,
         add_31_carry_3_, add_31_carry_4_, add_31_carry_5_, add_31_carry_6_,
         n22, n23, n24, n25, n26, n27, n28, n29, n30;

  add_4_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({in2[6:2], n23, n22}), .SUM(out3)
         );
  add_4_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, n29, temp2_2_, 
        temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_4_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, temp1_1_, temp1_0_}), .B({n26, in3[5:4], n25, n24, in3[1:0]}), .SUM(out2) );
  add_4_DW01_add_4 add_30 ( .A({in2[6:2], n23, n22}), .B({n26, in3[5:4], n25, 
        n24, in3[1:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}) );
  add_4_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX2 U1 ( .A(in2[0]), .Y(n22) );
  NAND2X8 U2 ( .A(add_31_n4), .B(add_31_n5), .Y(out[6]) );
  XOR2X1TH U3 ( .A(temp1_6_), .B(temp2_6_), .Y(add_31_n6) );
  ADDFXL U4 ( .A(temp1_5_), .B(temp2_5_), .CI(add_31_carry_5_), .CO(
        add_31_carry_6_), .S(out[5]) );
  BUFX2 U5 ( .A(in2[1]), .Y(n23) );
  BUFX2 U6 ( .A(in3[2]), .Y(n24) );
  INVX2TH U10 ( .A(add_31_carry_6_), .Y(n27) );
  BUFX2TH U14 ( .A(in3[3]), .Y(n25) );
  ADDFHXLTH U15 ( .A(temp1_4_), .B(temp2_4_), .CI(add_31_carry_4_), .CO(
        add_31_carry_5_), .S(out[4]) );
  NAND2X1 U16 ( .A(add_31_n6), .B(n27), .Y(add_31_n4) );
  ADDFHXLTH U17 ( .A(temp1_3_), .B(n29), .CI(add_31_carry_3_), .CO(
        add_31_carry_4_), .S(out[3]) );
  CLKBUFX1TH U18 ( .A(in3[6]), .Y(n26) );
  ADDFHXLTH U19 ( .A(temp1_2_), .B(temp2_2_), .CI(add_31_carry_2_), .CO(
        add_31_carry_3_), .S(out[2]) );
  CLKXOR2X1TH U20 ( .A(temp2_0_), .B(temp1_0_), .Y(out[0]) );
  INVXLTH U21 ( .A(add_31_n6), .Y(n28) );
  ADDFX1TH U22 ( .A(temp1_1_), .B(temp2_1_), .CI(add_31_n1), .CO(
        add_31_carry_2_), .S(out[1]) );
  AND2XLTH U23 ( .A(temp2_0_), .B(temp1_0_), .Y(add_31_n1) );
  CLKBUFX40 U13 ( .A(temp2_3_), .Y(n29) );
  AND2X8 U24 ( .A(n28), .B(add_31_carry_6_), .Y(n30) );
  CLKINVX40 U25 ( .A(n30), .Y(add_31_n5) );
endmodule


module tc_sm_19 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n25, n27, n28, n29, n30, n31, n32;

  BUFX18 U3 ( .A(in[6]), .Y(out[4]) );
  BUFX2TH U4 ( .A(in[6]), .Y(n25) );
  NOR3X1TH U5 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U6 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U7 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U8 ( .A(in[2]), .Y(n31) );
  XNOR2XLTH U9 ( .A(n31), .B(n11), .Y(n10) );
  NOR2XLTH U10 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U11 ( .A(n25), .Y(n27) );
  INVXLTH U12 ( .A(in[5]), .Y(n28) );
  INVXLTH U13 ( .A(in[4]), .Y(n29) );
  CLKINVX1TH U14 ( .A(in[3]), .Y(n30) );
  OAI33X4TH U16 ( .A0(in[4]), .A1(n25), .A2(in[5]), .B0(n13), .B1(n28), .B2(
        n29), .Y(n8) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n30), .B0(n25), .Y(n7) );
  OAI221XLTH U19 ( .A0(n27), .A1(n12), .B0(n25), .B1(n32), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U20 ( .A0(n27), .A1(n10), .B0(n25), .B1(n31), .C0(n8), .Y(out[2])
         );
  OAI211XLTH U21 ( .A0(n25), .A1(n30), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U22 ( .A0N(n30), .A1N(n9), .B0(n25), .Y(n13) );
endmodule


module tc_sm_18 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n19, n21, n22, n23, n24;

  OAI221XL U3 ( .A0(n21), .A1(n8), .B0(in[6]), .B1(n23), .C0(n6), .Y(out[2])
         );
  INVXL U4 ( .A(in[6]), .Y(n21) );
  OAI221XL U5 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n24), .C0(n6), .Y(out[1])
         );
  AOI21BX4 U6 ( .A0(in[6]), .A1(n11), .B0N(n19), .Y(n6) );
  NOR3X1TH U7 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  OAI2B11X2TH U8 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  OAI21BX4 U9 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n19) );
  INVXLTH U10 ( .A(in[2]), .Y(n23) );
  XOR2XLTH U11 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI211XLTH U13 ( .A0(in[6]), .A1(n22), .B0(n5), .C0(n6), .Y(out[3]) );
  OAI21XLTH U14 ( .A0(n7), .A1(n22), .B0(in[6]), .Y(n5) );
  XOR2XLTH U15 ( .A(in[0]), .B(n24), .Y(n10) );
  INVXLTH U16 ( .A(in[1]), .Y(n24) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  CLKBUFX1TH U18 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U19 ( .A(in[3]), .Y(n22) );
endmodule


module tc_sm_17 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n19, n21, n22, n23, n24, n25,
         n26;

  OA21XLTH U3 ( .A0(in[6]), .A1(n24), .B0(n7), .Y(n18) );
  NAND2XLTH U4 ( .A(n18), .B(n19), .Y(out[3]) );
  OAI2BB1X1 U5 ( .A0N(n24), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI221XL U6 ( .A0(n21), .A1(n12), .B0(in[6]), .B1(n26), .C0(n19), .Y(out[1])
         );
  INVXLTH U7 ( .A(in[6]), .Y(n21) );
  OAI221X1 U8 ( .A0(n21), .A1(n10), .B0(in[6]), .B1(n25), .C0(n19), .Y(out[2])
         );
  BUFX10 U9 ( .A(n8), .Y(n19) );
  INVXLTH U10 ( .A(in[4]), .Y(n23) );
  INVXLTH U11 ( .A(in[5]), .Y(n22) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n24) );
  NOR3X1TH U13 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  XNOR2XLTH U14 ( .A(n25), .B(n11), .Y(n10) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[2]), .Y(n25) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n19), .Y(out[0]) );
  INVXLTH U18 ( .A(in[1]), .Y(n26) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  CLKBUFX1TH U20 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U21 ( .A0(n9), .A1(n24), .B0(in[6]), .Y(n7) );
  OAI33X4 U22 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n22), .B2(
        n23), .Y(n8) );
endmodule


module tc_sm_16 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n22, n23, n24, n25, n27, n28,
         n29;

  INVX3TH U3 ( .A(in[4]), .Y(n22) );
  OAI221XL U4 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n8), .Y(out[1])
         );
  INVXL U5 ( .A(in[6]), .Y(n20) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  OAI211XLTH U10 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n8), .Y(out[3]) );
  INVXLTH U12 ( .A(in[5]), .Y(n21) );
  OAI21XLTH U13 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U14 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U16 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n12) );
  OAI221XLTH U18 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n8), .Y(
        out[2]) );
  XNOR2XLTH U19 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U21 ( .A(in[2]), .Y(n24) );
  AOI33X4 U6 ( .A0(n22), .A1(n28), .A2(n21), .B0(n29), .B1(in[5]), .B2(in[4]), 
        .Y(n27) );
  CLKINVX40 U7 ( .A(n27), .Y(n8) );
  CLKINVX40 U11 ( .A(in[6]), .Y(n28) );
  AOI21BX4 U22 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n29) );
endmodule


module total_3_test_43 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n56, w5_4_, n5, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_19 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_18 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_17 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_16 sm_tc_4 ( .out(in1), .in(in) );
  add_4 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), .in2(
        b1), .in3(c1), .in(in1) );
  tc_sm_19 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_18 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_17 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_16 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n45), .CK(clk), .RN(n5), 
        .Q(n56) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n41), .CK(clk), .RN(rst), 
        .Q(h) );
  SDFFRQX1TH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n42), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up2[2]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n42), .CK(clk), .RN(n5), 
        .Q(up3[3]) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQXLTH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n48), .CK(clk), .RN(n5), .Q(
        up1[0]) );
  SDFFRQX1TH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(up1[2]) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRQX1TH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n41), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRQX2 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up2[1]) );
  CLKBUFX4TH U3 ( .A(rst), .Y(n5) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n45), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  SDFFRHQX8 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n50), .CK(clk), .RN(rst), 
        .Q(up1[3]) );
  INVXLTH U36 ( .A(n44), .Y(n41) );
  INVXLTH U37 ( .A(n43), .Y(n42) );
  DLY1X1TH U38 ( .A(n47), .Y(n43) );
  DLY1X1TH U39 ( .A(n47), .Y(n44) );
  INVXLTH U40 ( .A(n44), .Y(n45) );
  INVXLTH U41 ( .A(n43), .Y(n46) );
  INVXLTH U42 ( .A(test_se), .Y(n47) );
  INVXLTH U43 ( .A(n44), .Y(n48) );
  INVXLTH U44 ( .A(n43), .Y(n49) );
  INVXLTH U45 ( .A(n44), .Y(n50) );
  INVXLTH U46 ( .A(n43), .Y(n51) );
  DLY1X1TH U47 ( .A(n56), .Y(up3[4]) );
endmodule


module sm_tc_15 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n32, n33, n36;

  NOR2X4 U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX3 U3 ( .A(in[4]), .Y(n32) );
  CLKBUFX1TH U4 ( .A(out[4]), .Y(out[6]) );
  XNOR2X2TH U5 ( .A(n36), .B(n8), .Y(n5) );
  NAND2XL U6 ( .A(n8), .B(n36), .Y(n7) );
  INVX1TH U7 ( .A(in[2]), .Y(n33) );
  OAI22X1 U8 ( .A0(in[4]), .A1(n36), .B0(n32), .B1(n5), .Y(out[2]) );
  CLKBUFX1TH U9 ( .A(in[0]), .Y(out[0]) );
  AOI31X2TH U10 ( .A0(n3), .A1(n4), .A2(n5), .B0(n32), .Y(out[4]) );
  AO21X1TH U11 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  OAI2BB2X4 U12 ( .B0(n32), .B1(n6), .A0N(in[1]), .A1N(n32), .Y(out[1]) );
  XNOR2X4 U13 ( .A(n7), .B(in[3]), .Y(n4) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2XLTH U16 ( .B0(n32), .B1(n4), .A0N(in[3]), .A1N(n32), .Y(out[3]) );
  CLKBUFX40 U17 ( .A(n33), .Y(n36) );
endmodule


module sm_tc_14 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n25, n29, n30, n33;

  XNOR2X1TH U2 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X2 U3 ( .B0(n30), .B1(n6), .A0N(in[1]), .A1N(n30), .Y(out[1]) );
  AO21X1 U5 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  BUFX2TH U6 ( .A(in[0]), .Y(out[0]) );
  NOR2X4 U7 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX4 U8 ( .A(in[2]), .Y(n29) );
  OAI2BB2X1 U9 ( .B0(n30), .B1(n4), .A0N(in[3]), .A1N(n30), .Y(out[3]) );
  INVX4 U10 ( .A(n25), .Y(n30) );
  BUFX6 U12 ( .A(in[4]), .Y(n25) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[6]) );
  NAND2XLTH U14 ( .A(n8), .B(n29), .Y(n7) );
  AOI31X2TH U15 ( .A0(n3), .A1(n4), .A2(n33), .B0(n30), .Y(out[4]) );
  CLKBUFX1TH U16 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U17 ( .AN(n6), .B(in[0]), .Y(n3) );
  OAI2B2X2 U4 ( .A1N(n25), .A0(n33), .B0(n25), .B1(n29), .Y(out[2]) );
  CLKBUFX40 U11 ( .A(n5), .Y(n33) );
  XNOR2X1 U18 ( .A(n29), .B(n8), .Y(n5) );
endmodule


module sm_tc_13 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n24, n25, n28, n29, n30, n31;

  XNOR2X1TH U3 ( .A(n7), .B(in[3]), .Y(n4) );
  XNOR2X1TH U4 ( .A(n25), .B(n8), .Y(n5) );
  OAI2BB2X4TH U5 ( .B0(n30), .B1(n6), .A0N(in[1]), .A1N(n30), .Y(out[1]) );
  INVX2 U6 ( .A(in[4]), .Y(n24) );
  AOI31X2 U7 ( .A0(n3), .A1(n4), .A2(n31), .B0(n30), .Y(out[4]) );
  OAI2BB2X2 U8 ( .B0(n30), .B1(n4), .A0N(in[3]), .A1N(n30), .Y(out[3]) );
  CLKBUFX1TH U9 ( .A(in[0]), .Y(out[0]) );
  NAND2XLTH U10 ( .A(n8), .B(n25), .Y(n7) );
  NOR2X4TH U11 ( .A(in[1]), .B(in[0]), .Y(n8) );
  INVX1TH U12 ( .A(in[2]), .Y(n25) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[5]) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[6]) );
  AO21XLTH U16 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKBUFX40 U2 ( .A(n24), .Y(n28) );
  OAI2B2X2 U17 ( .A1N(n29), .A0(n31), .B0(in[4]), .B1(n25), .Y(out[2]) );
  CLKINVX40 U18 ( .A(n28), .Y(n29) );
  CLKINVX40 U19 ( .A(n29), .Y(n30) );
  CLKBUFX40 U20 ( .A(n5), .Y(n31) );
endmodule


module sm_tc_12 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  OAI2BB2X2 U5 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  XNOR2X1 U2 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX1TH U3 ( .A(in[0]), .Y(out[0]) );
  CLKNAND2X2TH U4 ( .A(n8), .B(n21), .Y(n7) );
  INVXLTH U6 ( .A(out[4]), .Y(n18) );
  OAI22X1TH U7 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  NOR2X2TH U8 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U9 ( .A(n18), .Y(out[5]) );
  INVXLTH U10 ( .A(n18), .Y(out[6]) );
  OAI2BB2X1TH U11 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  CLKINVX1TH U12 ( .A(in[2]), .Y(n21) );
  CLKINVX2TH U13 ( .A(in[4]), .Y(n22) );
  AOI31X2TH U14 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U15 ( .AN(n6), .B(in[0]), .Y(n3) );
  XNOR2X1TH U16 ( .A(n21), .B(n8), .Y(n5) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_3_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_3_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_3_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(B[1]), .B(A[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR2X1TH U1 ( .A(B[6]), .B(A[6]), .Y(n2) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  CLKXOR2X12 U4 ( .A(n2), .B(carry[6]), .Y(SUM[6]) );
endmodule


module add_3_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n3;
  wire   [6:2] carry;

  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XNOR2X4TH U1 ( .A(n3), .B(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR2XLTH U3 ( .A(A[6]), .B(B[6]), .Y(n3) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_3_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4;
  wire   [6:2] carry;

  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  NAND3X4 U1 ( .A(n2), .B(n3), .C(n4), .Y(carry[2]) );
  NAND2X2 U2 ( .A(B[1]), .B(A[1]), .Y(n2) );
  NAND2X2TH U3 ( .A(B[1]), .B(n1), .Y(n3) );
  XOR3XL U4 ( .A(B[1]), .B(A[1]), .C(n1), .Y(SUM[1]) );
  NAND2X2 U5 ( .A(A[1]), .B(n1), .Y(n4) );
  AND2X1TH U6 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U7 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_3_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  XOR2X3TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_3 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n16, n17, n18, n19, n20;

  add_3_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n19, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in2[6:3], n16, n20, in2[0]}), .SUM(out3) );
  add_3_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_3_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n19, temp1_2_, 
        temp1_1_, temp1_0_}), .B({in3[6:3], n17, n18, in3[0]}), .SUM(out2) );
  add_3_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n19, temp1_2_, 
        temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_3_DW01_add_4 add_30 ( .A({in2[6:3], n16, n20, in2[0]}), .B({in3[6:3], 
        n17, n18, in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}) );
  add_3_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX2 U1 ( .A(in2[2]), .Y(n16) );
  BUFX6 U2 ( .A(in3[2]), .Y(n17) );
  CLKBUFX40 U3 ( .A(in3[1]), .Y(n18) );
  CLKBUFX40 U4 ( .A(temp1_3_), .Y(n19) );
  CLKBUFX40 U5 ( .A(in2[1]), .Y(n20) );
endmodule


module tc_sm_15 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31, n33;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(n33), .Y(n26) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(n33), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U11 ( .A(in[5]), .Y(n27) );
  INVXLTH U12 ( .A(in[4]), .Y(n28) );
  CLKINVX1TH U13 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U14 ( .A(n33), .Y(out[4]) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI21XLTH U16 ( .A0(n9), .A1(n29), .B0(n33), .Y(n7) );
  OAI221XLTH U17 ( .A0(n26), .A1(n12), .B0(n33), .B1(n31), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U18 ( .A0(n26), .A1(n10), .B0(n33), .B1(n30), .C0(n8), .Y(out[2])
         );
  OAI211XLTH U19 ( .A0(n33), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(n33), .Y(n13) );
  CLKBUFX40 U21 ( .A(in[6]), .Y(n33) );
endmodule


module tc_sm_14 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n25, n26, n27, n28, n29, n30, n31,
         n32, n34, n35, n36, n37, n39;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  NAND2X1TH U3 ( .A(n39), .B(n11), .Y(n25) );
  INVX5 U4 ( .A(n12), .Y(n26) );
  CLKAND2X8 U5 ( .A(n25), .B(n26), .Y(n6) );
  AOI2BB1X2 U6 ( .A0N(in[5]), .A1N(in[4]), .B0(n39), .Y(n12) );
  INVX2 U8 ( .A(n6), .Y(n29) );
  OAI211XLTH U9 ( .A0(n39), .A1(n35), .B0(n5), .C0(n6), .Y(out[3]) );
  NOR2X2 U10 ( .A(n34), .B(n10), .Y(n27) );
  OR3XLTH U11 ( .A(n27), .B(n28), .C(n29), .Y(out[1]) );
  OR3XLTH U12 ( .A(n30), .B(n31), .C(n32), .Y(out[2]) );
  NOR2X2 U13 ( .A(n8), .B(n34), .Y(n30) );
  OAI21XL U14 ( .A0(n7), .A1(n35), .B0(n39), .Y(n5) );
  NOR2XLTH U15 ( .A(n39), .B(n37), .Y(n28) );
  INVXLTH U16 ( .A(n39), .Y(n34) );
  NOR2XLTH U17 ( .A(n39), .B(n36), .Y(n31) );
  INVXLTH U18 ( .A(n6), .Y(n32) );
  XOR2X1TH U19 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR3X1TH U20 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U21 ( .A(n39), .Y(out[4]) );
  XOR2XLTH U22 ( .A(in[0]), .B(n37), .Y(n10) );
  INVXLTH U23 ( .A(in[1]), .Y(n37) );
  INVXLTH U24 ( .A(in[2]), .Y(n36) );
  NOR2XLTH U25 ( .A(in[0]), .B(in[1]), .Y(n9) );
  INVXLTH U26 ( .A(in[3]), .Y(n35) );
  NAND2BXLTH U27 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  CLKBUFX40 U28 ( .A(in[6]), .Y(n39) );
endmodule


module tc_sm_13 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n23, n24, n25, n26, n27, n28, n30, n31,
         n32;

  OAI211XL U3 ( .A0(in[6]), .A1(n26), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221XL U4 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n27), .C0(n8), .Y(out[2])
         );
  OAI221XL U5 ( .A0(n23), .A1(n12), .B0(in[6]), .B1(n28), .C0(n8), .Y(out[1])
         );
  CLKINVX1TH U7 ( .A(in[3]), .Y(n26) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVX2TH U9 ( .A(in[4]), .Y(n25) );
  INVXLTH U10 ( .A(in[1]), .Y(n28) );
  XNOR2XLTH U11 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U12 ( .A(n27), .B(n11), .Y(n10) );
  INVXLTH U13 ( .A(in[2]), .Y(n27) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n11) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI21XLTH U17 ( .A0(n9), .A1(n26), .B0(in[6]), .Y(n7) );
  INVXLTH U18 ( .A(in[6]), .Y(n23) );
  INVX2 U19 ( .A(in[5]), .Y(n24) );
  AOI33X4 U6 ( .A0(n25), .A1(n31), .A2(n24), .B0(n32), .B1(in[4]), .B2(in[5]), 
        .Y(n30) );
  CLKINVX40 U20 ( .A(n30), .Y(n8) );
  CLKINVX40 U21 ( .A(in[6]), .Y(n31) );
  AOI21BX4 U22 ( .A0(n26), .A1(n9), .B0N(in[6]), .Y(n32) );
endmodule


module tc_sm_12 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n21, n23, n24, n25, n26;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  CLKINVX1TH U3 ( .A(in[6]), .Y(n23) );
  OAI211XLTH U4 ( .A0(in[6]), .A1(n24), .B0(n5), .C0(n6), .Y(out[3]) );
  AOI21BX4 U5 ( .A0(in[6]), .A1(n11), .B0N(n21), .Y(n6) );
  OAI21BX2 U6 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n21) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n9) );
  XOR2XLTH U10 ( .A(in[0]), .B(n26), .Y(n10) );
  INVXLTH U11 ( .A(in[1]), .Y(n26) );
  OAI21XLTH U12 ( .A0(n7), .A1(n24), .B0(in[6]), .Y(n5) );
  INVXLTH U13 ( .A(in[3]), .Y(n24) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  OAI221XLTH U16 ( .A0(n23), .A1(n8), .B0(in[6]), .B1(n25), .C0(n6), .Y(out[2]) );
  INVXLTH U17 ( .A(in[2]), .Y(n25) );
  XOR2XLTH U18 ( .A(in[2]), .B(n9), .Y(n8) );
  OAI221XLTH U19 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n26), .C0(n6), .Y(
        out[1]) );
endmodule


module total_3_test_44 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n6, n7, n46, n47, n48, n49, n50, n51, n52, n53, n54, n56;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_15 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_14 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_13 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_12 sm_tc_4 ( .out(in1), .in(in) );
  add_3 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), .in2(
        b1), .in3(c1), .in(in1) );
  tc_sm_15 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_14 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_13 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_12 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up3[0]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n53), .CK(clk), .RN(n7), 
        .Q(up3[3]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up2[3]) );
  SDFFRQXLTH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up2[1]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up2[0]) );
  SDFFRQXLTH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n47), .CK(clk), .RN(n6), 
        .Q(up2[2]) );
  SDFFRQXLTH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n47), .CK(clk), .RN(n6), .Q(
        up1[0]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(up3[2]) );
  SDFFRQXL up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(up1[2]) );
  SDFFRQX2 up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n52), .CK(clk), .RN(n6), 
        .Q(up2[4]) );
  SDFFRQX2 up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n53), .CK(clk), .RN(n6), 
        .Q(up3[4]) );
  SDFFRQX4 up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up1[4]) );
  SDFFRQX1 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n49), .CK(clk), .RN(n7), 
        .Q(up1[3]) );
  CLKBUFX1TH U3 ( .A(rst), .Y(n7) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n6) );
  SDFFRX4 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n50), .CK(clk), .RN(n6), 
        .Q(n54) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up3[1]) );
  SDFFRX4 h_reg ( .D(w5_4_), .SI(test_si), .SE(n52), .CK(clk), .RN(n7), .Q(h)
         );
  DLY1X1TH U37 ( .A(n51), .Y(n46) );
  INVXLTH U38 ( .A(n46), .Y(n47) );
  INVXLTH U39 ( .A(n46), .Y(n48) );
  DLY1X1TH U40 ( .A(test_se), .Y(n49) );
  DLY1X1TH U41 ( .A(test_se), .Y(n50) );
  INVXLTH U42 ( .A(test_se), .Y(n51) );
  INVXLTH U43 ( .A(n46), .Y(n52) );
  INVXLTH U44 ( .A(n46), .Y(n53) );
  CLKINVX40 U45 ( .A(n54), .Y(n56) );
  CLKINVX40 U46 ( .A(n56), .Y(up1[1]) );
endmodule


module sm_tc_11 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n23, n26, n27, n28, n29, n30;

  OAI22X1 U11 ( .A0(in[4]), .A1(n23), .B0(n22), .B1(n28), .Y(out[2]) );
  XNOR2X2TH U2 ( .A(n7), .B(in[3]), .Y(n4) );
  AOI31X1 U3 ( .A0(n3), .A1(n28), .A2(n4), .B0(n22), .Y(out[4]) );
  OAI2BB2X4 U4 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  INVX4 U5 ( .A(in[4]), .Y(n22) );
  NOR2X4 U6 ( .A(in[1]), .B(n26), .Y(n8) );
  CLKBUFX1TH U7 ( .A(n26), .Y(out[0]) );
  INVX2 U9 ( .A(in[2]), .Y(n23) );
  CLKBUFX1TH U10 ( .A(out[4]), .Y(out[6]) );
  NOR2BXLTH U13 ( .AN(n6), .B(n26), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  NAND2XLTH U15 ( .A(n8), .B(n23), .Y(n7) );
  XOR2X1 U8 ( .A(n23), .B(n30), .Y(n5) );
  CLKBUFX40 U12 ( .A(in[0]), .Y(n26) );
  AO2B2BX4 U16 ( .A0(n27), .A1N(n4), .B0(in[3]), .B1N(n27), .Y(out[3]) );
  CLKINVX40 U17 ( .A(n22), .Y(n27) );
  CLKBUFX40 U18 ( .A(n5), .Y(n28) );
  AOI21BX4 U19 ( .A0(n26), .A1(in[1]), .B0N(n30), .Y(n29) );
  CLKINVX40 U20 ( .A(n29), .Y(n6) );
  CLKINVX40 U21 ( .A(n8), .Y(n30) );
endmodule


module sm_tc_10 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n39, n3, n4, n5, n6, n8, n25, n29, n30, n33, n34, n36, n37, n38;

  XNOR2X1 U2 ( .A(n30), .B(n8), .Y(n5) );
  NOR2X3 U4 ( .A(in[1]), .B(in[0]), .Y(n8) );
  BUFX6 U5 ( .A(n5), .Y(n25) );
  AOI31X2TH U7 ( .A0(n3), .A1(n4), .A2(n25), .B0(n37), .Y(n39) );
  INVX1TH U8 ( .A(in[2]), .Y(n30) );
  CLKBUFX1TH U9 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2X1TH U10 ( .B0(n37), .B1(n4), .A0N(in[3]), .A1N(n37), .Y(out[3]) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  OAI22X1TH U12 ( .A0(n36), .A1(n30), .B0(n37), .B1(n25), .Y(out[2]) );
  CLKBUFX1TH U13 ( .A(in[0]), .Y(out[0]) );
  NOR2BXLTH U14 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVX2TH U15 ( .A(in[4]), .Y(n29) );
  OAI2BB2X2 U16 ( .B0(n37), .B1(n6), .A0N(in[1]), .A1N(n37), .Y(out[1]) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKBUFX40 U3 ( .A(n29), .Y(n33) );
  CLKINVX40 U6 ( .A(n39), .Y(n34) );
  CLKINVX40 U18 ( .A(n34), .Y(out[4]) );
  CLKINVX40 U19 ( .A(n33), .Y(n36) );
  CLKINVX40 U20 ( .A(n36), .Y(n37) );
  XOR2X1 U21 ( .A(n38), .B(in[3]), .Y(n4) );
  CLKAND2X12 U22 ( .A(n8), .B(n30), .Y(n38) );
endmodule


module sm_tc_9 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n27, n31, n32, n35, n36;

  BUFX2 U2 ( .A(in[1]), .Y(n27) );
  XNOR2X2TH U4 ( .A(n31), .B(n8), .Y(n5) );
  OAI2BB2X1TH U5 ( .B0(n32), .B1(n4), .A0N(in[3]), .A1N(n32), .Y(out[3]) );
  CLKBUFX1TH U6 ( .A(in[0]), .Y(out[0]) );
  AOI31X2TH U7 ( .A0(n3), .A1(n4), .A2(n5), .B0(n32), .Y(out[4]) );
  XNOR2X2TH U8 ( .A(n7), .B(in[3]), .Y(n4) );
  INVX2TH U9 ( .A(in[4]), .Y(n32) );
  NOR2BXLTH U10 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U12 ( .A(out[4]), .Y(out[6]) );
  NAND2XLTH U13 ( .A(n8), .B(n31), .Y(n7) );
  CLKINVX1TH U14 ( .A(in[2]), .Y(n31) );
  OAI2BB2X2 U15 ( .B0(n32), .B1(n6), .A0N(n27), .A1N(n32), .Y(out[1]) );
  OAI22XL U17 ( .A0(in[4]), .A1(n31), .B0(n32), .B1(n5), .Y(out[2]) );
  AOI21BX4 U3 ( .A0(in[0]), .A1(n27), .B0N(n36), .Y(n35) );
  CLKINVX40 U16 ( .A(n35), .Y(n6) );
  OR2X8 U18 ( .A(n27), .B(in[0]), .Y(n36) );
  CLKINVX40 U19 ( .A(n36), .Y(n8) );
endmodule


module sm_tc_8 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n22, n25, n26;

  OAI2BB2X2 U5 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n26), .Y(out[1]) );
  NOR2BX1 U9 ( .AN(n6), .B(in[0]), .Y(n3) );
  NAND2X2TH U2 ( .A(n8), .B(n25), .Y(n7) );
  XNOR2X1 U3 ( .A(n7), .B(in[3]), .Y(n4) );
  AOI31X2 U4 ( .A0(n3), .A1(n4), .A2(n5), .B0(n26), .Y(out[4]) );
  XNOR2X1 U6 ( .A(n25), .B(n8), .Y(n5) );
  CLKBUFX1TH U7 ( .A(in[0]), .Y(out[0]) );
  NOR2X2TH U8 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI2BB2X1TH U10 ( .B0(n26), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  INVXLTH U11 ( .A(n22), .Y(out[5]) );
  OAI22X1TH U12 ( .A0(in[4]), .A1(n25), .B0(n26), .B1(n5), .Y(out[2]) );
  CLKINVX2TH U13 ( .A(in[4]), .Y(n26) );
  INVXLTH U14 ( .A(out[4]), .Y(n22) );
  CLKINVX1TH U15 ( .A(in[2]), .Y(n25) );
  INVXLTH U16 ( .A(n22), .Y(out[6]) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_2_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1TH U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_2_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n3, n4, n5, n6, n7;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n5), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR2XLTH U4 ( .A(B[4]), .B(A[4]), .Y(n1) );
  XOR2X1TH U5 ( .A(n1), .B(carry[4]), .Y(SUM[4]) );
  AND2XLTH U6 ( .A(B[0]), .B(A[0]), .Y(n5) );
  CLKXOR2X1TH U7 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2XLTH U8 ( .A(A[4]), .B(B[4]), .Y(n4) );
  AND2X8 U1 ( .A(carry[4]), .B(B[4]), .Y(n6) );
  CLKINVX40 U2 ( .A(n6), .Y(n3) );
  AND2X8 U3 ( .A(carry[4]), .B(A[4]), .Y(n7) );
  NAND3BX4 U9 ( .AN(n7), .B(n3), .C(n4), .Y(carry[5]) );
endmodule


module add_2_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_2_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_2_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n5, n1, n3, n4;
  wire   [6:2] carry;

  ADDFHX2TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(n5) );
  XOR3XLTH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX2 U1_4 ( .A(carry[4]), .B(B[4]), .CI(A[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKBUFX40 U1 ( .A(n5), .Y(SUM[5]) );
  DLY1X1TH U3 ( .A(n4), .Y(n3) );
  XNOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(n4) );
  CLKINVX40 U5 ( .A(n3), .Y(SUM[0]) );
endmodule


module add_2_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X1TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX2TH U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_2 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;

  add_2_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, n30, temp1_2_, 
        temp1_1_, n27}), .B({in2[6], n25, in2[4], n29, in2[2], n26, in2[0]}), 
        .SUM(out3) );
  add_2_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, n28, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_2_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, n30, temp1_2_, 
        temp1_1_, n27}), .B({in3[6:5], n21, in3[3], n23, n20, n24}), .SUM(out2) );
  add_2_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, n30, temp1_2_, 
        temp1_1_, n27}), .B({temp2_6_, temp2_5_, n28, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .SUM(out) );
  add_2_DW01_add_4 add_30 ( .A({in2[6], n25, in2[4], n29, in2[2], n26, in2[0]}), .B({in3[6:5], n21, in3[3], n23, n20, n24}), .SUM({temp2_6_, temp2_5_, 
        temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_}) );
  add_2_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  BUFX10 U1 ( .A(in3[1]), .Y(n20) );
  CLKBUFX1TH U2 ( .A(in3[4]), .Y(n21) );
  INVX2 U3 ( .A(in3[2]), .Y(n22) );
  INVX2 U4 ( .A(n22), .Y(n23) );
  CLKBUFX40 U5 ( .A(in3[0]), .Y(n24) );
  CLKBUFX40 U6 ( .A(in2[5]), .Y(n25) );
  CLKBUFX40 U13 ( .A(in2[1]), .Y(n26) );
  CLKBUFX40 U14 ( .A(temp1_0_), .Y(n27) );
  CLKBUFX40 U15 ( .A(temp2_4_), .Y(n28) );
  CLKBUFX40 U16 ( .A(in2[3]), .Y(n29) );
  CLKBUFX40 U17 ( .A(temp1_3_), .Y(n30) );
endmodule


module tc_sm_11 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n25, n27, n28, n29, n30, n31, n32;

  CLKBUFX2TH U3 ( .A(in[6]), .Y(n25) );
  NOR3X1TH U4 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U5 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U6 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U7 ( .A(in[2]), .Y(n31) );
  XNOR2XLTH U8 ( .A(n31), .B(n11), .Y(n10) );
  NOR2XLTH U9 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U10 ( .A(n25), .Y(n27) );
  OAI33X4TH U11 ( .A0(in[4]), .A1(n25), .A2(in[5]), .B0(n13), .B1(n28), .B2(
        n29), .Y(n8) );
  INVXLTH U12 ( .A(in[5]), .Y(n28) );
  INVXLTH U13 ( .A(in[4]), .Y(n29) );
  CLKINVX1TH U14 ( .A(in[3]), .Y(n30) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U16 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI221XLTH U17 ( .A0(n27), .A1(n12), .B0(n25), .B1(n32), .C0(n8), .Y(out[1])
         );
  OAI221XLTH U18 ( .A0(n27), .A1(n10), .B0(n25), .B1(n31), .C0(n8), .Y(out[2])
         );
  OAI21XLTH U19 ( .A0(n9), .A1(n30), .B0(n25), .Y(n7) );
  OAI211XLTH U20 ( .A0(n25), .A1(n30), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U21 ( .A0N(n30), .A1N(n9), .B0(n25), .Y(n13) );
endmodule


module tc_sm_10 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n10, n11, n12, n27, n28, n29, n30, n31, n32, n34, n35, n36,
         n37, n38, n39, n40;

  BUFX2 U3 ( .A(n34), .Y(out[4]) );
  OAI211X2TH U4 ( .A0(out[4]), .A1(n30), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221X2 U8 ( .A0(n27), .A1(n10), .B0(out[4]), .B1(n31), .C0(n8), .Y(out[2])
         );
  OAI221X2TH U10 ( .A0(n27), .A1(n12), .B0(out[4]), .B1(n32), .C0(n8), .Y(
        out[1]) );
  INVX1TH U11 ( .A(in[5]), .Y(n28) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n30) );
  XNOR2XLTH U14 ( .A(n31), .B(n11), .Y(n10) );
  NAND2BXLTH U15 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U16 ( .A(in[2]), .Y(n31) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U18 ( .A(in[1]), .Y(n32) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVX2 U20 ( .A(in[4]), .Y(n29) );
  INVXLTH U21 ( .A(n34), .Y(n27) );
  CLKBUFX40 U5 ( .A(in[6]), .Y(n34) );
  OR3XLTH U6 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n35) );
  INVXLTH U7 ( .A(n35), .Y(n36) );
  OAI21BX4 U9 ( .A0(n36), .A1(n30), .B0N(n38), .Y(n7) );
  AOI33X4 U13 ( .A0(n29), .A1(n38), .A2(n28), .B0(n40), .B1(in[5]), .B2(n39), 
        .Y(n37) );
  CLKINVX40 U22 ( .A(n37), .Y(n8) );
  CLKINVX40 U23 ( .A(n34), .Y(n38) );
  CLKINVX40 U24 ( .A(n29), .Y(n39) );
  AOI21BX4 U25 ( .A0(n30), .A1(n36), .B0N(in[6]), .Y(n40) );
endmodule


module tc_sm_9 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n34, n35, n36, n37, n39, n40,
         n41;

  CLKINVX4TH U3 ( .A(in[6]), .Y(n34) );
  AOI21X1 U4 ( .A0(n5), .A1(n35), .B0(n6), .Y(out[3]) );
  NOR4X1 U5 ( .A(n7), .B(n34), .C(n8), .D(n35), .Y(n6) );
  NAND2XLTH U7 ( .A(n35), .B(n7), .Y(n13) );
  AOI2BB1X4 U9 ( .A0N(in[6]), .A1N(n5), .B0(n8), .Y(n10) );
  CLKINVX1TH U10 ( .A(in[3]), .Y(n35) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U12 ( .A(in[6]), .Y(out[4]) );
  XOR2XLTH U13 ( .A(in[0]), .B(n37), .Y(n12) );
  INVXLTH U14 ( .A(in[1]), .Y(n37) );
  INVXLTH U15 ( .A(in[2]), .Y(n36) );
  XOR2XLTH U16 ( .A(in[2]), .B(n11), .Y(n9) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI221XLTH U18 ( .A0(n34), .A1(n12), .B0(in[6]), .B1(n37), .C0(n10), .Y(
        out[1]) );
  OAI221XLTH U19 ( .A0(n34), .A1(n9), .B0(in[6]), .B1(n36), .C0(n10), .Y(
        out[2]) );
  NAND2BXLTH U20 ( .AN(in[0]), .B(n10), .Y(out[0]) );
  DLY1X1TH U6 ( .A(in[4]), .Y(n39) );
  OR3X8 U8 ( .A(in[5]), .B(in[6]), .C(n39), .Y(n40) );
  CLKINVX40 U21 ( .A(n40), .Y(n5) );
  AND3X8 U22 ( .A(in[5]), .B(n13), .C(n39), .Y(n41) );
  NOR2X8 U23 ( .A(n41), .B(n34), .Y(n8) );
endmodule


module tc_sm_8 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n23, n25, n26, n27, n28, n30;

  OAI2B11X2 U7 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  AOI21BX4 U3 ( .A0(in[6]), .A1(n11), .B0N(n23), .Y(n6) );
  INVXLTH U4 ( .A(in[6]), .Y(n25) );
  NOR3X1TH U5 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  CLKBUFX1TH U6 ( .A(in[6]), .Y(out[4]) );
  OAI21XLTH U8 ( .A0(n7), .A1(n26), .B0(in[6]), .Y(n5) );
  INVXLTH U9 ( .A(in[3]), .Y(n26) );
  XOR2XLTH U10 ( .A(in[0]), .B(n28), .Y(n10) );
  INVXLTH U11 ( .A(in[1]), .Y(n28) );
  INVXLTH U12 ( .A(in[2]), .Y(n27) );
  XOR2XLTH U13 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U14 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI21BX1 U15 ( .A0(in[5]), .A1(in[4]), .B0N(in[6]), .Y(n23) );
  OAI221XLTH U16 ( .A0(n25), .A1(n10), .B0(in[6]), .B1(n28), .C0(n6), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n30), .A1(n8), .B0(in[6]), .B1(n27), .C0(n6), .Y(out[2]) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n26), .B0(n5), .C0(n6), .Y(out[3]) );
  INVXLTH U20 ( .A(in[6]), .Y(n30) );
endmodule


module total_3_test_45 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n65, n66, w5_4_, n4, n5, n6, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n60;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_11 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_10 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_9 sm_tc_3 ( .out(c1), .in({c[4:1], n4}) );
  sm_tc_8 sm_tc_4 ( .out(in1), .in(in) );
  add_2 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), .in2(
        b1), .in3(c1), .in(in1) );
  tc_sm_11 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_10 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_9 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_8 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n52), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  SDFFRQXLTH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n54), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n55), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up1[2]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n47), .CK(clk), .RN(n6), 
        .Q(n66) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n47), .CK(clk), .RN(n5), 
        .Q(up1[3]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n54), .CK(clk), .RN(n5), .Q(
        up1[0]) );
  SDFFRQX1TH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n57), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  SDFFRQX2TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n48), .CK(clk), .RN(n6), 
        .Q(n65) );
  SDFFRQX2TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n52), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n56), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  BUFX2 U3 ( .A(c[0]), .Y(n4) );
  CLKBUFX1TH U4 ( .A(rst), .Y(n6) );
  CLKBUFX4TH U5 ( .A(rst), .Y(n5) );
  SDFFRX4 up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n57), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n55), .CK(clk), .RN(n5), 
        .Q(up2[1]) );
  SDFFRX4 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n56), .CK(clk), .RN(n5), 
        .Q(up2[2]) );
  SDFFRX4 up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n51), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRX4 h_reg ( .D(w5_4_), .SI(test_si), .SE(n51), .CK(clk), .RN(n6), .Q(h)
         );
  INVXLTH U38 ( .A(n50), .Y(n47) );
  INVXLTH U39 ( .A(n49), .Y(n48) );
  DLY1X1TH U40 ( .A(n53), .Y(n49) );
  DLY1X1TH U41 ( .A(n53), .Y(n50) );
  INVXLTH U42 ( .A(n50), .Y(n51) );
  INVXLTH U43 ( .A(n49), .Y(n52) );
  INVXLTH U44 ( .A(test_se), .Y(n53) );
  INVXLTH U45 ( .A(n50), .Y(n54) );
  INVXLTH U46 ( .A(n49), .Y(n55) );
  INVXLTH U47 ( .A(n50), .Y(n56) );
  INVXLTH U48 ( .A(n49), .Y(n57) );
  CLKINVX40 U49 ( .A(n65), .Y(n60) );
  CLKINVX40 U50 ( .A(n60), .Y(up3[4]) );
  DLY1X1TH U51 ( .A(n66), .Y(up3[3]) );
endmodule


module sm_tc_7 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n28, n29, n32, n33, n34;

  OAI2BB2X2 U5 ( .B0(n28), .B1(n6), .A0N(n33), .A1N(n28), .Y(out[1]) );
  XNOR2X1 U2 ( .A(n29), .B(n8), .Y(n5) );
  NOR2X6 U3 ( .A(n33), .B(in[0]), .Y(n8) );
  INVX4 U4 ( .A(in[4]), .Y(n28) );
  CLKBUFX1TH U7 ( .A(in[0]), .Y(out[0]) );
  AO21X4TH U8 ( .A0(in[0]), .A1(n33), .B0(n8), .Y(n6) );
  INVX1TH U9 ( .A(n32), .Y(n29) );
  OAI2BB2XLTH U10 ( .B0(n4), .B1(n28), .A0N(in[3]), .A1N(n28), .Y(out[3]) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  AOI31X2TH U12 ( .A0(n3), .A1(n4), .A2(n5), .B0(n28), .Y(out[4]) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX40 U6 ( .A(in[2]), .Y(n32) );
  OAI2BB2X2 U15 ( .B0(n28), .B1(n5), .A0N(n28), .A1N(n32), .Y(out[2]) );
  CLKBUFX40 U16 ( .A(in[1]), .Y(n33) );
  XOR2X1 U17 ( .A(n34), .B(in[3]), .Y(n4) );
  CLKAND2X12 U18 ( .A(n29), .B(n8), .Y(n34) );
endmodule


module sm_tc_6 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n17, n18, n19, n23, n24;

  XNOR2X2 U2 ( .A(n24), .B(n8), .Y(n5) );
  CLKBUFX2TH U3 ( .A(in[4]), .Y(n17) );
  XNOR2X2 U4 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKBUFX2TH U5 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X2TH U6 ( .B0(n23), .B1(n6), .A0N(in[1]), .A1N(n23), .Y(out[1]) );
  CLKAND2X2TH U7 ( .A(n18), .B(n19), .Y(out[5]) );
  NAND3X2TH U8 ( .A(n3), .B(n4), .C(n5), .Y(n18) );
  AO21X2 U9 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  NOR2X4 U10 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI22X1TH U11 ( .A0(n24), .A1(n17), .B0(n23), .B1(n5), .Y(out[2]) );
  NAND2XLTH U12 ( .A(n8), .B(n24), .Y(n7) );
  INVX2 U13 ( .A(in[2]), .Y(n24) );
  BUFX2TH U14 ( .A(out[5]), .Y(out[4]) );
  INVXLTH U15 ( .A(n23), .Y(n19) );
  CLKBUFX1TH U16 ( .A(out[5]), .Y(out[6]) );
  INVX6 U17 ( .A(n17), .Y(n23) );
  OAI2BB2X1TH U18 ( .B0(n23), .B1(n4), .A0N(in[3]), .A1N(n23), .Y(out[3]) );
  NOR2BXLTH U19 ( .AN(n6), .B(in[0]), .Y(n3) );
endmodule


module sm_tc_5 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n21, n22, n23, n27, n28;

  INVX4TH U2 ( .A(n23), .Y(n27) );
  OR2XLTH U3 ( .A(n23), .B(n28), .Y(n21) );
  OR2X2 U4 ( .A(n27), .B(n5), .Y(n22) );
  NAND2X2 U5 ( .A(n21), .B(n22), .Y(out[2]) );
  BUFX2 U6 ( .A(in[4]), .Y(n23) );
  INVX2 U7 ( .A(in[2]), .Y(n28) );
  XNOR2X1TH U8 ( .A(n28), .B(n8), .Y(n5) );
  NOR2X6 U9 ( .A(in[1]), .B(in[0]), .Y(n8) );
  AOI31X2 U10 ( .A0(n3), .A1(n4), .A2(n5), .B0(n27), .Y(out[4]) );
  OAI2BB2X1 U11 ( .B0(n27), .B1(n4), .A0N(in[3]), .A1N(n27), .Y(out[3]) );
  XNOR2X1TH U12 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X4 U13 ( .B0(n27), .B1(n6), .A0N(in[1]), .A1N(n27), .Y(out[1]) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[6]) );
  NAND2XL U15 ( .A(n8), .B(n28), .Y(n7) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U17 ( .A(out[4]), .Y(out[5]) );
  BUFX2TH U18 ( .A(in[0]), .Y(out[0]) );
  AO21XLTH U19 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module sm_tc_4 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  NOR2X2 U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  NAND2XL U3 ( .A(n8), .B(n21), .Y(n7) );
  AOI31X2TH U4 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  XNOR2X1 U5 ( .A(n21), .B(n8), .Y(n5) );
  OAI2BB2X2TH U6 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  OAI22X1TH U7 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  CLKBUFX1TH U8 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X2TH U9 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKINVX2TH U10 ( .A(in[4]), .Y(n22) );
  INVXLTH U11 ( .A(n18), .Y(out[6]) );
  CLKINVX1TH U12 ( .A(in[2]), .Y(n21) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U14 ( .A(out[4]), .Y(n18) );
  INVXLTH U15 ( .A(n18), .Y(out[5]) );
  XNOR2X1TH U16 ( .A(n7), .B(in[3]), .Y(n4) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_1_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_1_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n4, n1, n2;
  wire   [6:2] carry;

  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n4) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKINVX40 U3 ( .A(n4), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_1_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module add_1_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, n1;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry_2_), .S(SUM[1]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry_6_), .Y(SUM[6]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_1_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7;
  wire   [6:2] carry;

  CLKXOR2X1TH U3 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CLKXOR2X2TH U1 ( .A(n1), .B(carry[6]), .Y(SUM[6]) );
  XOR2XLTH U2 ( .A(B[6]), .B(A[6]), .Y(n1) );
  AND2XLTH U4 ( .A(B[0]), .B(A[0]), .Y(n2) );
  CLKBUFX40 U5 ( .A(n4), .Y(n3) );
  DLY1X1TH U6 ( .A(n2), .Y(n4) );
  XOR3X4 U7 ( .A(A[1]), .B(B[1]), .C(n3), .Y(SUM[1]) );
  NAND2X8 U8 ( .A(A[1]), .B(B[1]), .Y(n5) );
  NAND2X8 U9 ( .A(A[1]), .B(n3), .Y(n6) );
  NAND2X8 U10 ( .A(B[1]), .B(n3), .Y(n7) );
  NAND3X8 U11 ( .A(n5), .B(n6), .C(n7), .Y(carry[2]) );
endmodule


module add_1_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  XOR3X2 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_1 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n17, n18, n19, n20, n21, n22, n23, n24;

  add_1_DW01_add_0 add_34 ( .A({temp1_6_, n22, temp1_4_, temp1_3_, n23, 
        temp1_1_, temp1_0_}), .B({in2[6:3], n20, n24, in2[0]}), .SUM(out3) );
  add_1_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .B({in[6:3], n18, n17, in[0]}), .SUM(
        out1) );
  add_1_DW01_add_2 add_32 ( .A({temp1_6_, n22, temp1_4_, temp1_3_, n23, 
        temp1_1_, temp1_0_}), .B({in3[6:2], n21, in3[0]}), .SUM(out2) );
  add_1_DW01_add_3 add_31 ( .A({temp1_6_, n22, temp1_4_, temp1_3_, n23, 
        temp1_1_, temp1_0_}), .B({temp2_6_, temp2_5_, temp2_4_, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_1_DW01_add_4 add_30 ( .A({in2[6:3], n20, n24, in2[0]}), .B({in3[6:2], 
        n21, in3[0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_1_DW01_add_5 add_29 ( .A({in[6:2], n17, in[0]}), .B(in1), .SUM({temp1_6_, 
        temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  INVX2 U1 ( .A(in2[2]), .Y(n19) );
  BUFX2TH U2 ( .A(in[1]), .Y(n17) );
  CLKBUFX1TH U3 ( .A(in[2]), .Y(n18) );
  INVX2TH U4 ( .A(n19), .Y(n20) );
  BUFX4 U5 ( .A(in3[1]), .Y(n21) );
  CLKBUFX40 U6 ( .A(temp1_5_), .Y(n22) );
  CLKBUFX40 U13 ( .A(temp1_2_), .Y(n23) );
  CLKBUFX40 U14 ( .A(in2[1]), .Y(n24) );
endmodule


module tc_sm_7 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n24, n25, n26, n27, n28, n29;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n28) );
  XNOR2XLTH U7 ( .A(n28), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U9 ( .A(in[6]), .Y(n24) );
  OAI33X4TH U10 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n25), .B2(
        n26), .Y(n8) );
  INVXLTH U11 ( .A(in[4]), .Y(n26) );
  INVXLTH U12 ( .A(in[5]), .Y(n25) );
  OAI21XLTH U13 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  CLKINVX1TH U14 ( .A(in[3]), .Y(n27) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  OAI221XLTH U16 ( .A0(n24), .A1(n12), .B0(in[6]), .B1(n29), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(
        out[2]) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n27), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_6 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n34, n35, n36, n38, n39;

  OAI221XL U3 ( .A0(n34), .A1(n12), .B0(in[6]), .B1(n36), .C0(n11), .Y(out[1])
         );
  OAI31X2TH U4 ( .A0(n34), .A1(n8), .A2(n10), .B0(n11), .Y(n9) );
  AO21XL U5 ( .A0(n34), .A1(in[2]), .B0(n9), .Y(out[2]) );
  CLKNAND2X2TH U6 ( .A(n4), .B(n5), .Y(out[3]) );
  OAI31X1 U7 ( .A0(n7), .A1(n8), .A2(n35), .B0(in[6]), .Y(n4) );
  NAND3X6 U8 ( .A(in[5]), .B(in[4]), .C(n13), .Y(n7) );
  INVX16 U9 ( .A(in[6]), .Y(n34) );
  CLKNAND2X8 U10 ( .A(n6), .B(n7), .Y(n11) );
  OR3X2 U11 ( .A(in[5]), .B(in[6]), .C(in[4]), .Y(n6) );
  INVX2TH U13 ( .A(in[3]), .Y(n35) );
  NOR3X4TH U14 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n8) );
  XOR2XLTH U15 ( .A(in[0]), .B(n36), .Y(n12) );
  INVXLTH U16 ( .A(in[1]), .Y(n36) );
  OA21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(in[2]), .Y(n10) );
  CLKBUFX1TH U18 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U19 ( .AN(in[0]), .B(n11), .Y(out[0]) );
  OA21X4 U12 ( .A0(in[3]), .A1(n6), .B0(n34), .Y(n38) );
  CLKINVX40 U20 ( .A(n38), .Y(n5) );
  AOI21BX4 U21 ( .A0(n8), .A1(n35), .B0N(n39), .Y(n13) );
  CLKINVX40 U22 ( .A(n34), .Y(n39) );
endmodule


module tc_sm_5 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n18, n20, n21, n22, n23, n24, n25;

  OAI211XL U3 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n18), .Y(out[3]) );
  OAI2BB1X4 U4 ( .A0N(n23), .A1N(n9), .B0(in[6]), .Y(n13) );
  OAI221XL U5 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n18), .Y(out[2])
         );
  BUFX8 U6 ( .A(n8), .Y(n18) );
  OAI221XL U7 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n18), .Y(out[1])
         );
  INVXLTH U8 ( .A(in[6]), .Y(n20) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U10 ( .A(in[3]), .Y(n23) );
  OAI21XLTH U11 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  INVXLTH U12 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n12) );
  XNOR2XLTH U14 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U15 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U16 ( .A(in[2]), .Y(n24) );
  CLKBUFX1TH U17 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U18 ( .AN(in[0]), .B(n18), .Y(out[0]) );
  OAI33X4 U19 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n21), .B2(
        n22), .Y(n8) );
  INVXL U20 ( .A(in[5]), .Y(n21) );
  INVXL U21 ( .A(in[4]), .Y(n22) );
endmodule


module tc_sm_4 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n19, n21, n22, n23, n24, n26, n27, n28,
         n29;

  OAI221XL U4 ( .A0(n19), .A1(n12), .B0(in[6]), .B1(n24), .C0(n8), .Y(out[1])
         );
  OAI221XL U5 ( .A0(n19), .A1(n10), .B0(in[6]), .B1(n23), .C0(n8), .Y(out[2])
         );
  OAI211XL U6 ( .A0(in[6]), .A1(n22), .B0(n7), .C0(n8), .Y(out[3]) );
  NOR3X1TH U7 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n22) );
  INVXLTH U9 ( .A(in[6]), .Y(n19) );
  CLKBUFX1TH U10 ( .A(in[6]), .Y(out[4]) );
  XNOR2XLTH U11 ( .A(n23), .B(n11), .Y(n10) );
  NOR2XLTH U12 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U13 ( .A(in[2]), .Y(n23) );
  OAI21XLTH U14 ( .A0(n9), .A1(n22), .B0(in[6]), .Y(n7) );
  INVXLTH U15 ( .A(in[1]), .Y(n24) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXL U20 ( .A(in[4]), .Y(n21) );
  AOI33X4 U3 ( .A0(n21), .A1(n27), .A2(n28), .B0(n29), .B1(in[5]), .B2(in[4]), 
        .Y(n26) );
  CLKINVX40 U18 ( .A(n26), .Y(n8) );
  CLKINVX40 U19 ( .A(in[6]), .Y(n27) );
  CLKINVX40 U21 ( .A(in[5]), .Y(n28) );
  AOI21BX4 U22 ( .A0(n22), .A1(n9), .B0N(in[6]), .Y(n29) );
endmodule


module total_3_test_46 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   w5_4_, n6, n7, n8, n43, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_7 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_6 sm_tc_2 ( .out(b1), .in({b[4:2], n43, b[0]}) );
  sm_tc_5 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_4 sm_tc_4 ( .out(in1), .in(in) );
  add_1 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), .in2(
        b1), .in3({c1[6:3], n6, c1[1:0]}), .in(in1) );
  tc_sm_7 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_6 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_5 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_4 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n51), .CK(clk), .RN(n7), 
        .Q(up3[0]) );
  SDFFRQX1TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n58), .CK(clk), .RN(n7), 
        .Q(up1[4]) );
  SDFFRHQX1TH up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n55), .CK(clk), .RN(n7), 
        .Q(up1[1]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(h), .SE(n57), .CK(clk), .RN(n7), .Q(
        up1[0]) );
  SDFFRQX1TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n50), .CK(clk), .RN(n7), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n58), .CK(clk), .RN(n8), 
        .Q(up3[3]) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n57), .CK(clk), .RN(n7), 
        .Q(up2[3]) );
  SDFFRQXLTH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n50), .CK(clk), .RN(n8), 
        .Q(up3[4]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n55), .CK(clk), .RN(n7), 
        .Q(up3[1]) );
  SDFFRQXLTH up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n50), .CK(clk), .RN(n7), 
        .Q(up3[2]) );
  CLKBUFX1TH U3 ( .A(c1[2]), .Y(n6) );
  CLKBUFX4TH U4 ( .A(rst), .Y(n7) );
  CLKBUFX1TH U5 ( .A(rst), .Y(n8) );
  SDFFRX4 up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n55), .CK(clk), .RN(n7), 
        .Q(up2[0]) );
  SDFFRX4 up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n51), .CK(clk), .RN(n7), 
        .Q(up2[1]) );
  SDFFRHQX8 up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n59), .CK(clk), .RN(n7), 
        .Q(up1[3]) );
  SDFFRX4 h_reg ( .D(w5_4_), .SI(test_si), .SE(n55), .CK(clk), .RN(n8), .Q(h)
         );
  SDFFRX4 up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n51), .CK(clk), .RN(n7), 
        .Q(up2[2]) );
  SDFFRHQX8 up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n59), .CK(clk), .RN(n7), 
        .Q(up1[2]) );
  CLKBUFX40 U38 ( .A(b[1]), .Y(n43) );
  DLY1X1TH U39 ( .A(n53), .Y(n50) );
  DLY1X1TH U40 ( .A(n54), .Y(n51) );
  DLY1X1TH U41 ( .A(n56), .Y(n52) );
  INVXLTH U42 ( .A(n52), .Y(n53) );
  INVXLTH U43 ( .A(n56), .Y(n54) );
  DLY1X1TH U44 ( .A(test_se), .Y(n55) );
  INVXLTH U45 ( .A(test_se), .Y(n56) );
  INVXLTH U46 ( .A(n52), .Y(n57) );
  INVXLTH U47 ( .A(n52), .Y(n58) );
  INVXLTH U48 ( .A(n52), .Y(n59) );
endmodule


module sm_tc_3 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n8, n22, n26, n27, n30, n31;

  BUFX2 U2 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X2 U3 ( .B0(n26), .B1(n6), .A0N(in[1]), .A1N(n31), .Y(out[1]) );
  OAI22X1 U4 ( .A0(n22), .A1(n27), .B0(n26), .B1(n5), .Y(out[2]) );
  INVX4 U5 ( .A(n22), .Y(n26) );
  BUFX10 U6 ( .A(in[4]), .Y(n22) );
  AOI31X1 U8 ( .A0(n3), .A1(n5), .A2(n4), .B0(n31), .Y(out[4]) );
  XNOR2X2TH U9 ( .A(n27), .B(n8), .Y(n5) );
  NOR2X6TH U10 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKBUFX1TH U11 ( .A(out[4]), .Y(out[6]) );
  INVX2TH U12 ( .A(in[2]), .Y(n27) );
  AO21X4 U13 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  OAI2BB2XLTH U15 ( .B0(n31), .B1(n4), .A0N(in[3]), .A1N(n26), .Y(out[3]) );
  NOR2BXLTH U16 ( .AN(n6), .B(in[0]), .Y(n3) );
  XOR2X1 U7 ( .A(n30), .B(in[3]), .Y(n4) );
  CLKAND2X12 U17 ( .A(n8), .B(n27), .Y(n30) );
  INVX4 U18 ( .A(n22), .Y(n31) );
endmodule


module sm_tc_2 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n23, n24, n27, n28, n29, n30;

  NOR2BXLTH U2 ( .AN(n6), .B(in[0]), .Y(n3) );
  XNOR2X2 U3 ( .A(n24), .B(n8), .Y(n5) );
  INVX3 U4 ( .A(in[4]), .Y(n23) );
  NOR2X3 U5 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKNAND2X2TH U6 ( .A(n8), .B(n24), .Y(n7) );
  XNOR2X2TH U8 ( .A(n7), .B(in[3]), .Y(n4) );
  CLKINVX1TH U9 ( .A(in[2]), .Y(n24) );
  OAI2BB2X4TH U10 ( .B0(n28), .B1(n6), .A0N(n29), .A1N(n28), .Y(out[1]) );
  CLKBUFX1TH U11 ( .A(in[0]), .Y(out[0]) );
  OAI2BB2X1TH U12 ( .B0(n28), .B1(n4), .A0N(in[3]), .A1N(n28), .Y(out[3]) );
  CLKBUFX1TH U13 ( .A(out[4]), .Y(out[6]) );
  BUFX2TH U14 ( .A(out[4]), .Y(out[5]) );
  AOI31X4 U16 ( .A0(n3), .A1(n4), .A2(n5), .B0(n28), .Y(out[4]) );
  OAI2BB2X2 U7 ( .B0(n28), .B1(n5), .A0N(n23), .A1N(in[2]), .Y(out[2]) );
  CLKINVX40 U15 ( .A(n23), .Y(n27) );
  CLKINVX40 U17 ( .A(n27), .Y(n28) );
  DLY1X1TH U18 ( .A(in[1]), .Y(n29) );
  AOI21X8 U19 ( .A0(in[0]), .A1(n29), .B0(n8), .Y(n30) );
  CLKINVX40 U20 ( .A(n30), .Y(n6) );
endmodule


module sm_tc_1 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n28, n32, n33, n36, n37, n38;

  OAI2BB2X2 U3 ( .B0(n38), .B1(n4), .A0N(in[3]), .A1N(n38), .Y(out[3]) );
  INVX2 U2 ( .A(in[2]), .Y(n33) );
  XNOR2X1TH U4 ( .A(n7), .B(in[3]), .Y(n4) );
  OAI2BB2X4 U5 ( .B0(n38), .B1(n6), .A0N(n36), .A1N(n38), .Y(out[1]) );
  NOR2X2 U6 ( .A(n36), .B(in[0]), .Y(n8) );
  XNOR2X1 U7 ( .A(n33), .B(n8), .Y(n5) );
  BUFX2TH U8 ( .A(in[0]), .Y(out[0]) );
  AO21X4 U9 ( .A0(in[0]), .A1(n36), .B0(n8), .Y(n6) );
  INVXLTH U10 ( .A(n38), .Y(n28) );
  INVX2TH U11 ( .A(in[4]), .Y(n32) );
  CLKNAND2X2 U12 ( .A(n8), .B(n33), .Y(n7) );
  NOR2BXLTH U13 ( .AN(n6), .B(in[0]), .Y(n3) );
  CLKBUFX1TH U14 ( .A(out[4]), .Y(out[5]) );
  CLKBUFX1TH U15 ( .A(out[4]), .Y(out[6]) );
  OAI22X4 U16 ( .A0(n28), .A1(n33), .B0(n38), .B1(n5), .Y(out[2]) );
  AOI31X4 U17 ( .A0(n3), .A1(n4), .A2(n5), .B0(n38), .Y(out[4]) );
  CLKBUFX40 U18 ( .A(in[1]), .Y(n36) );
  CLKINVX40 U19 ( .A(n32), .Y(n37) );
  CLKINVX40 U20 ( .A(n37), .Y(n38) );
endmodule


module sm_tc_0 ( out, in );
  output [6:0] out;
  input [4:0] in;
  wire   n3, n4, n5, n6, n7, n8, n18, n21, n22;

  NOR2X4TH U2 ( .A(in[1]), .B(in[0]), .Y(n8) );
  OAI22X1TH U3 ( .A0(in[4]), .A1(n21), .B0(n22), .B1(n5), .Y(out[2]) );
  OAI2BB2X1TH U4 ( .B0(n22), .B1(n6), .A0N(in[1]), .A1N(n22), .Y(out[1]) );
  CLKBUFX1TH U5 ( .A(in[0]), .Y(out[0]) );
  INVXLTH U6 ( .A(n18), .Y(out[6]) );
  NAND2XLTH U7 ( .A(n8), .B(n21), .Y(n7) );
  CLKINVX2TH U8 ( .A(in[4]), .Y(n22) );
  CLKINVX1TH U9 ( .A(in[2]), .Y(n21) );
  AOI31X2TH U10 ( .A0(n3), .A1(n4), .A2(n5), .B0(n22), .Y(out[4]) );
  NOR2BXLTH U11 ( .AN(n6), .B(in[0]), .Y(n3) );
  INVXLTH U12 ( .A(n18), .Y(out[5]) );
  INVXLTH U13 ( .A(out[4]), .Y(n18) );
  OAI2BB2X1TH U14 ( .B0(n22), .B1(n4), .A0N(in[3]), .A1N(n22), .Y(out[3]) );
  XNOR2X1TH U15 ( .A(n21), .B(n8), .Y(n5) );
  XNOR2X1TH U16 ( .A(n7), .B(in[3]), .Y(n4) );
  AO21XLTH U17 ( .A0(in[0]), .A1(in[1]), .B0(n8), .Y(n6) );
endmodule


module add_0_DW01_add_0 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X4TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_0_DW01_add_1 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  CLKXOR2X2TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CLKAND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_0_DW01_add_2 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(n1), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  AND2XLTH U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1TH U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module add_0_DW01_add_3 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2;
  wire   [6:2] carry;

  ADDFX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHXLTH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFHXLTH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHXLTH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFHXLTH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CLKXOR2X1TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR3X2 U3 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(n2) );
  CLKINVX40 U4 ( .A(n2), .Y(SUM[6]) );
endmodule


module add_0_DW01_add_4 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n1, n2, n4, n5, n6, n7, n8, n9;
  wire   [6:2] carry;

  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFHX1TH U1_1 ( .A(n1), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2TH U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFHX2TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X3 U2 ( .A(n2), .B(carry[4]), .Y(SUM[4]) );
  AND2X4TH U7 ( .A(A[0]), .B(B[0]), .Y(n1) );
  NAND2XLTH U8 ( .A(A[4]), .B(B[4]), .Y(n5) );
  AND2X8 U3 ( .A(carry[4]), .B(B[4]), .Y(n6) );
  CLKINVX40 U4 ( .A(n6), .Y(n4) );
  XOR2X1 U5 ( .A(n7), .B(n8), .Y(n2) );
  CLKINVX40 U6 ( .A(B[4]), .Y(n7) );
  CLKINVX40 U9 ( .A(A[4]), .Y(n8) );
  NAND3BX4 U10 ( .AN(n9), .B(n4), .C(n5), .Y(carry[5]) );
  CLKAND2X12 U11 ( .A(carry[4]), .B(A[4]), .Y(n9) );
endmodule


module add_0_DW01_add_5 ( A, B, SUM );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  wire   n3, n1;
  wire   [6:2] carry;

  ADDFX1TH U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1TH U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1TH U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(n3) );
  XOR3X2TH U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .Y(SUM[6]) );
  ADDFHX1TH U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CLKXOR2X2TH U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2XLTH U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKBUFX40 U3 ( .A(n3), .Y(SUM[2]) );
endmodule


module add_0 ( out1, out2, out3, out, in1, in2, in3, in );
  output [6:0] out1;
  output [6:0] out2;
  output [6:0] out3;
  output [6:0] out;
  input [6:0] in1;
  input [6:0] in2;
  input [6:0] in3;
  input [6:0] in;
  wire   temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, temp2_1_, temp2_0_,
         temp1_6_, temp1_5_, temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_,
         n22, n23, n24, n25;

  add_0_DW01_add_0 add_34 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n25, temp1_0_}), .B({in2[6:4], n23, in2[2:0]}), .SUM(out3)
         );
  add_0_DW01_add_1 add_33 ( .A({temp2_6_, temp2_5_, n22, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}), .B(in), .SUM(out1) );
  add_0_DW01_add_2 add_32 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n25, temp1_0_}), .B({in3[6:4], n24, in3[2:0]}), .SUM(out2)
         );
  add_0_DW01_add_3 add_31 ( .A({temp1_6_, temp1_5_, temp1_4_, temp1_3_, 
        temp1_2_, n25, temp1_0_}), .B({temp2_6_, temp2_5_, n22, temp2_3_, 
        temp2_2_, temp2_1_, temp2_0_}), .SUM(out) );
  add_0_DW01_add_4 add_30 ( .A({in2[6:4], n23, in2[2:0]}), .B({in3[6:4], n24, 
        in3[2:0]}), .SUM({temp2_6_, temp2_5_, temp2_4_, temp2_3_, temp2_2_, 
        temp2_1_, temp2_0_}) );
  add_0_DW01_add_5 add_29 ( .A(in), .B(in1), .SUM({temp1_6_, temp1_5_, 
        temp1_4_, temp1_3_, temp1_2_, temp1_1_, temp1_0_}) );
  CLKBUFX2 U1 ( .A(temp2_4_), .Y(n22) );
  CLKBUFX40 U2 ( .A(in2[3]), .Y(n23) );
  CLKBUFX40 U3 ( .A(in3[3]), .Y(n24) );
  CLKBUFX40 U4 ( .A(temp1_1_), .Y(n25) );
endmodule


module tc_sm_3 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n13, n26, n27, n28, n29, n30, n31;

  NOR3X1TH U3 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U4 ( .A(in[1]), .Y(n31) );
  XNOR2XLTH U5 ( .A(in[0]), .B(in[1]), .Y(n12) );
  INVXLTH U6 ( .A(in[2]), .Y(n30) );
  XNOR2XLTH U7 ( .A(n30), .B(n11), .Y(n10) );
  NOR2XLTH U8 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI33X4TH U9 ( .A0(in[4]), .A1(in[6]), .A2(in[5]), .B0(n13), .B1(n27), .B2(
        n28), .Y(n8) );
  INVXLTH U10 ( .A(in[5]), .Y(n27) );
  INVXLTH U11 ( .A(in[4]), .Y(n28) );
  CLKINVX1TH U12 ( .A(in[3]), .Y(n29) );
  CLKBUFX1TH U13 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U14 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  INVXLTH U15 ( .A(in[6]), .Y(n26) );
  OAI221XLTH U16 ( .A0(n26), .A1(n12), .B0(in[6]), .B1(n31), .C0(n8), .Y(
        out[1]) );
  OAI221XLTH U17 ( .A0(n26), .A1(n10), .B0(in[6]), .B1(n30), .C0(n8), .Y(
        out[2]) );
  OAI21XLTH U18 ( .A0(n9), .A1(n29), .B0(in[6]), .Y(n7) );
  OAI211XLTH U19 ( .A0(in[6]), .A1(n29), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI2BB1XLTH U20 ( .A0N(n29), .A1N(n9), .B0(in[6]), .Y(n13) );
endmodule


module tc_sm_2 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n8, n9, n10, n11, n12, n20, n21, n23, n24, n25, n26, n27, n28,
         n29, n31, n32, n33;

  NAND2BX2 U3 ( .AN(in[0]), .B(n8), .Y(out[0]) );
  OAI211X2 U4 ( .A0(in[6]), .A1(n27), .B0(n7), .C0(n8), .Y(out[3]) );
  OAI221X2 U5 ( .A0(n24), .A1(n10), .B0(in[6]), .B1(n28), .C0(n8), .Y(out[2])
         );
  NAND3XL U6 ( .A(n20), .B(n21), .C(n8), .Y(out[1]) );
  OR2XLTH U7 ( .A(n24), .B(n12), .Y(n20) );
  OR2XLTH U8 ( .A(in[6]), .B(n29), .Y(n21) );
  INVXLTH U9 ( .A(in[6]), .Y(n24) );
  NOR3X1TH U11 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  INVXLTH U12 ( .A(n9), .Y(n23) );
  XNOR2XLTH U13 ( .A(n28), .B(n11), .Y(n10) );
  OAI21XLTH U14 ( .A0(n9), .A1(n27), .B0(in[6]), .Y(n7) );
  CLKBUFX1TH U15 ( .A(in[6]), .Y(out[4]) );
  INVX2 U16 ( .A(in[5]), .Y(n25) );
  INVXLTH U17 ( .A(in[3]), .Y(n27) );
  INVXLTH U18 ( .A(in[1]), .Y(n29) );
  XNOR2XLTH U19 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NOR2XLTH U20 ( .A(in[0]), .B(in[1]), .Y(n11) );
  INVXLTH U21 ( .A(in[2]), .Y(n28) );
  INVXL U23 ( .A(in[4]), .Y(n26) );
  AOI33X4 U10 ( .A0(n26), .A1(n32), .A2(n25), .B0(n33), .B1(in[5]), .B2(in[4]), 
        .Y(n31) );
  CLKINVX40 U22 ( .A(n31), .Y(n8) );
  CLKINVX40 U24 ( .A(in[6]), .Y(n32) );
  OA21X4 U25 ( .A0(in[3]), .A1(n23), .B0(in[6]), .Y(n33) );
endmodule


module tc_sm_1 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n7, n9, n10, n11, n12, n20, n21, n22, n23, n24, n25, n27, n28, n29,
         n30;

  OAI211X2 U3 ( .A0(in[6]), .A1(n23), .B0(n7), .C0(n30), .Y(out[3]) );
  OAI221X1 U5 ( .A0(n20), .A1(n12), .B0(in[6]), .B1(n25), .C0(n30), .Y(out[1])
         );
  OAI221X1 U6 ( .A0(n20), .A1(n10), .B0(in[6]), .B1(n24), .C0(n30), .Y(out[2])
         );
  INVXLTH U7 ( .A(in[6]), .Y(n20) );
  CLKINVX1TH U8 ( .A(in[3]), .Y(n23) );
  NOR3X1TH U9 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n9) );
  CLKBUFX1TH U10 ( .A(in[6]), .Y(out[4]) );
  INVXLTH U11 ( .A(in[1]), .Y(n25) );
  XNOR2XLTH U12 ( .A(n24), .B(n11), .Y(n10) );
  NOR2XLTH U13 ( .A(in[0]), .B(in[1]), .Y(n11) );
  OAI21XLTH U14 ( .A0(n9), .A1(n23), .B0(in[6]), .Y(n7) );
  INVXLTH U15 ( .A(in[2]), .Y(n24) );
  XNOR2XLTH U16 ( .A(in[0]), .B(in[1]), .Y(n12) );
  NAND2BXLTH U17 ( .AN(in[0]), .B(n30), .Y(out[0]) );
  INVXL U19 ( .A(in[5]), .Y(n21) );
  INVXL U20 ( .A(in[4]), .Y(n22) );
  AOI33X4 U4 ( .A0(n22), .A1(n28), .A2(n21), .B0(n29), .B1(in[5]), .B2(in[4]), 
        .Y(n27) );
  CLKINVX40 U18 ( .A(in[6]), .Y(n28) );
  AOI21BX4 U21 ( .A0(n23), .A1(n9), .B0N(in[6]), .Y(n29) );
  CLKINVX40 U22 ( .A(n27), .Y(n30) );
endmodule


module tc_sm_0 ( out, in );
  output [4:0] out;
  input [6:0] in;
  wire   n5, n6, n7, n8, n9, n10, n11, n20, n21, n23, n24, n25, n26, n28, n29;

  NAND2X1 U3 ( .A(in[6]), .B(n11), .Y(n21) );
  OAI221XL U4 ( .A0(n23), .A1(n10), .B0(in[6]), .B1(n26), .C0(n6), .Y(out[1])
         );
  AND2X6TH U5 ( .A(n21), .B(n20), .Y(n6) );
  INVXLTH U7 ( .A(in[6]), .Y(n23) );
  NOR3X1TH U8 ( .A(in[1]), .B(in[2]), .C(in[0]), .Y(n7) );
  OAI2B11XLTH U9 ( .A1N(n7), .A0(in[3]), .B0(in[4]), .C0(in[5]), .Y(n11) );
  CLKBUFX1TH U10 ( .A(in[6]), .Y(out[4]) );
  NAND2BXLTH U11 ( .AN(in[0]), .B(n6), .Y(out[0]) );
  XOR2XLTH U12 ( .A(in[0]), .B(n26), .Y(n10) );
  INVXLTH U13 ( .A(in[1]), .Y(n26) );
  OAI221XLTH U14 ( .A0(n23), .A1(n8), .B0(in[6]), .B1(n25), .C0(n6), .Y(out[2]) );
  INVXLTH U15 ( .A(in[2]), .Y(n25) );
  XOR2XLTH U16 ( .A(in[2]), .B(n9), .Y(n8) );
  NOR2XLTH U17 ( .A(in[0]), .B(in[1]), .Y(n9) );
  OAI21XLTH U19 ( .A0(n7), .A1(n24), .B0(in[6]), .Y(n5) );
  INVXLTH U20 ( .A(in[3]), .Y(n24) );
  OAI2B11X4 U6 ( .A1N(n28), .A0(n24), .B0(n5), .C0(n6), .Y(out[3]) );
  CLKINVX40 U18 ( .A(in[6]), .Y(n28) );
  AOI2BB1X4 U21 ( .A0N(in[5]), .A1N(in[4]), .B0(in[6]), .Y(n29) );
  CLKINVX40 U22 ( .A(n29), .Y(n20) );
endmodule


module total_3_test_47 ( h, up1, up2, up3, clk, rst, a, b, c, in, test_si, 
        test_se );
  output [4:0] up1;
  output [4:0] up2;
  output [4:0] up3;
  input [4:0] a;
  input [4:0] b;
  input [4:0] c;
  input [4:0] in;
  input clk, rst, test_si, test_se;
  output h;
  wire   n59, n60, n61, w5_4_, n4, n5, n6, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n53, n55, n57;
  wire   [6:0] a1;
  wire   [6:0] b1;
  wire   [6:0] c1;
  wire   [6:0] in1;
  wire   [6:0] w66;
  wire   [6:0] w77;
  wire   [6:0] w88;
  wire   [6:0] w55;
  wire   [4:0] w6;
  wire   [4:0] w7;
  wire   [4:0] w8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  sm_tc_3 sm_tc_1 ( .out(a1), .in(a) );
  sm_tc_2 sm_tc_2 ( .out(b1), .in(b) );
  sm_tc_1 sm_tc_3 ( .out(c1), .in(c) );
  sm_tc_0 sm_tc_4 ( .out(in1), .in(in) );
  add_0 add_1 ( .out1(w66), .out2(w77), .out3(w88), .out(w55), .in1(a1), .in2(
        b1), .in3({c1[6:1], n4}), .in(in1) );
  tc_sm_3 tc_sm_1 ( .out({w5_4_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}), .in(w55) );
  tc_sm_2 tc_sm_2 ( .out(w6), .in(w66) );
  tc_sm_1 tc_sm_3 ( .out(w7), .in(w77) );
  tc_sm_0 tc_sm_4 ( .out(w8), .in(w88) );
  SDFFRQXLTH up2_reg_3_ ( .D(w7[3]), .SI(up2[2]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up2[3]) );
  SDFFRQXLTH up2_reg_1_ ( .D(w7[1]), .SI(up2[0]), .SE(n42), .CK(clk), .RN(n5), 
        .Q(up2[1]) );
  SDFFRQX1TH up1_reg_0_ ( .D(w6[0]), .SI(n57), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up1[0]) );
  SDFFRQXLTH h_reg ( .D(w5_4_), .SI(test_si), .SE(n45), .CK(clk), .RN(n6), .Q(
        n59) );
  SDFFRQXLTH up2_reg_0_ ( .D(w7[0]), .SI(up1[4]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up2[0]) );
  SDFFRQX2TH up3_reg_4_ ( .D(w8[4]), .SI(up3[3]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(n60) );
  SDFFRQXLTH up3_reg_3_ ( .D(w8[3]), .SI(up3[2]), .SE(n44), .CK(clk), .RN(n5), 
        .Q(n61) );
  SDFFRQX2TH up1_reg_4_ ( .D(w6[4]), .SI(up1[3]), .SE(n49), .CK(clk), .RN(n5), 
        .Q(up1[4]) );
  SDFFRQX1TH up2_reg_2_ ( .D(w7[2]), .SI(up2[1]), .SE(n48), .CK(clk), .RN(n5), 
        .Q(up2[2]) );
  SDFFRQXLTH up3_reg_1_ ( .D(w8[1]), .SI(up3[0]), .SE(n50), .CK(clk), .RN(n5), 
        .Q(up3[1]) );
  SDFFRQXLTH up1_reg_3_ ( .D(w6[3]), .SI(up1[2]), .SE(n49), .CK(clk), .RN(n6), 
        .Q(up1[3]) );
  SDFFRQXLTH up1_reg_2_ ( .D(w6[2]), .SI(up1[1]), .SE(n46), .CK(clk), .RN(n6), 
        .Q(up1[2]) );
  SDFFRQX1TH up2_reg_4_ ( .D(w7[4]), .SI(up2[3]), .SE(n42), .CK(clk), .RN(n5), 
        .Q(up2[4]) );
  SDFFRQXLTH up3_reg_0_ ( .D(w8[0]), .SI(up2[4]), .SE(n45), .CK(clk), .RN(n5), 
        .Q(up3[0]) );
  SDFFRHQX2 up1_reg_1_ ( .D(w6[1]), .SI(up1[0]), .SE(n46), .CK(clk), .RN(n5), 
        .Q(up1[1]) );
  CLKBUFX2TH U3 ( .A(c1[0]), .Y(n4) );
  CLKBUFX1TH U4 ( .A(rst), .Y(n6) );
  CLKBUFX4TH U5 ( .A(rst), .Y(n5) );
  SDFFRX4 up3_reg_2_ ( .D(w8[2]), .SI(up3[1]), .SE(n44), .CK(clk), .RN(n5), 
        .Q(up3[2]) );
  DLY1X1TH U38 ( .A(n43), .Y(n41) );
  INVXLTH U39 ( .A(n43), .Y(n42) );
  DLY1X1TH U40 ( .A(n47), .Y(n43) );
  INVXLTH U41 ( .A(n43), .Y(n44) );
  INVXLTH U42 ( .A(n47), .Y(n45) );
  DLY1X1TH U43 ( .A(test_se), .Y(n46) );
  INVXLTH U44 ( .A(test_se), .Y(n47) );
  INVXLTH U45 ( .A(n41), .Y(n48) );
  INVXLTH U46 ( .A(n41), .Y(n49) );
  INVXLTH U47 ( .A(n43), .Y(n50) );
  CLKINVX40 U48 ( .A(n60), .Y(n53) );
  CLKINVX40 U49 ( .A(n53), .Y(up3[4]) );
  INVXLTH U50 ( .A(n59), .Y(n55) );
  INVXLTH U51 ( .A(n55), .Y(h) );
  INVXLTH U52 ( .A(n55), .Y(n57) );
  DLY1X1TH U53 ( .A(n61), .Y(up3[3]) );
endmodule


module iteration_test_1 ( h1, h2, h3, h4, h5, h6, h7, h8, h9, h10, h11, h12, 
        h13, h14, h15, h16, h17, h18, h19, h20, h21, h22, h23, h24, h25, h26, 
        h27, h28, h29, h30, h31, h32, h33, h34, h35, h36, h37, h38, h39, h40, 
        h41, h42, h43, h44, h45, h46, h47, h48, clk, rst, i1, i2, i3, i4, i5, 
        i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20, 
        i21, i22, i23, i24, i25, i26, i27, i28, i29, i30, i31, i32, i33, i34, 
        i35, i36, i37, i38, i39, i40, i41, i42, i43, i44, i45, i46, i47, i48, 
        test_si, test_so, test_se );
  input [4:0] i1;
  input [4:0] i2;
  input [4:0] i3;
  input [4:0] i4;
  input [4:0] i5;
  input [4:0] i6;
  input [4:0] i7;
  input [4:0] i8;
  input [4:0] i9;
  input [4:0] i10;
  input [4:0] i11;
  input [4:0] i12;
  input [4:0] i13;
  input [4:0] i14;
  input [4:0] i15;
  input [4:0] i16;
  input [4:0] i17;
  input [4:0] i18;
  input [4:0] i19;
  input [4:0] i20;
  input [4:0] i21;
  input [4:0] i22;
  input [4:0] i23;
  input [4:0] i24;
  input [4:0] i25;
  input [4:0] i26;
  input [4:0] i27;
  input [4:0] i28;
  input [4:0] i29;
  input [4:0] i30;
  input [4:0] i31;
  input [4:0] i32;
  input [4:0] i33;
  input [4:0] i34;
  input [4:0] i35;
  input [4:0] i36;
  input [4:0] i37;
  input [4:0] i38;
  input [4:0] i39;
  input [4:0] i40;
  input [4:0] i41;
  input [4:0] i42;
  input [4:0] i43;
  input [4:0] i44;
  input [4:0] i45;
  input [4:0] i46;
  input [4:0] i47;
  input [4:0] i48;
  input clk, rst, test_si, test_se;
  output h1, h2, h3, h4, h5, h6, h7, h8, h9, h10, h11, h12, h13, h14, h15, h16,
         h17, h18, h19, h20, h21, h22, h23, h24, h25, h26, h27, h28, h29, h30,
         h31, h32, h33, h34, h35, h36, h37, h38, h39, h40, h41, h42, h43, h44,
         h45, h46, h47, h48, test_so;
  wire   up48_3_3_, up48_3_2_, up48_3_1_, up48_3_0_, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120;
  wire   [4:0] c1_1;
  wire   [4:0] c1_2;
  wire   [4:0] c1_3;
  wire   [4:0] c1_4;
  wire   [4:0] c1_5;
  wire   [4:0] c1_6;
  wire   [4:0] up3_1;
  wire   [4:0] up6_1;
  wire   [4:0] up18_1;
  wire   [4:0] up20_1;
  wire   [4:0] up26_1;
  wire   [4:0] up27_1;
  wire   [4:0] c2_1;
  wire   [4:0] c2_2;
  wire   [4:0] c2_3;
  wire   [4:0] c2_4;
  wire   [4:0] c2_5;
  wire   [4:0] c2_6;
  wire   [4:0] up4_1;
  wire   [4:0] up5_1;
  wire   [4:0] up17_1;
  wire   [4:0] up19_1;
  wire   [4:0] up25_1;
  wire   [4:0] up28_1;
  wire   [4:0] c3_1;
  wire   [4:0] c3_2;
  wire   [4:0] c3_3;
  wire   [4:0] c3_4;
  wire   [4:0] c3_5;
  wire   [4:0] c3_6;
  wire   [4:0] up4_2;
  wire   [4:0] up14_1;
  wire   [4:0] up16_1;
  wire   [4:0] up27_2;
  wire   [4:0] up29_1;
  wire   [4:0] up31_1;
  wire   [4:0] c4_1;
  wire   [4:0] c4_2;
  wire   [4:0] c4_3;
  wire   [4:0] c4_4;
  wire   [4:0] c4_5;
  wire   [4:0] c4_6;
  wire   [4:0] up3_2;
  wire   [4:0] up13_1;
  wire   [4:0] up15_1;
  wire   [4:0] up28_2;
  wire   [4:0] up30_1;
  wire   [4:0] up32_1;
  wire   [4:0] c5_1;
  wire   [4:0] c5_2;
  wire   [4:0] c5_3;
  wire   [4:0] c5_4;
  wire   [4:0] c5_5;
  wire   [4:0] c5_6;
  wire   [4:0] up7_1;
  wire   [4:0] up9_1;
  wire   [4:0] up12_1;
  wire   [4:0] up29_2;
  wire   [4:0] up31_2;
  wire   [4:0] up33_1;
  wire   [4:0] c6_1;
  wire   [4:0] c6_2;
  wire   [4:0] c6_3;
  wire   [4:0] c6_4;
  wire   [4:0] c6_5;
  wire   [4:0] c6_6;
  wire   [4:0] up8_1;
  wire   [4:0] up10_1;
  wire   [4:0] up11_1;
  wire   [4:0] up30_2;
  wire   [4:0] up32_2;
  wire   [4:0] up34_1;
  wire   [4:0] c7_1;
  wire   [4:0] c7_2;
  wire   [4:0] c7_3;
  wire   [4:0] c7_4;
  wire   [4:0] c7_5;
  wire   [4:0] c7_6;
  wire   [4:0] up2_1;
  wire   [4:0] up6_2;
  wire   [4:0] up18_2;
  wire   [4:0] up20_2;
  wire   [4:0] up29_3;
  wire   [4:0] up31_3;
  wire   [4:0] c8_1;
  wire   [4:0] c8_2;
  wire   [4:0] c8_3;
  wire   [4:0] c8_4;
  wire   [4:0] c8_5;
  wire   [4:0] c8_6;
  wire   [4:0] up1_1;
  wire   [4:0] up5_2;
  wire   [4:0] up17_2;
  wire   [4:0] up19_2;
  wire   [4:0] up30_3;
  wire   [4:0] up32_3;
  wire   [4:0] c9_1;
  wire   [4:0] c9_2;
  wire   [4:0] c9_3;
  wire   [4:0] c9_4;
  wire   [4:0] c9_5;
  wire   [4:0] c9_6;
  wire   [4:0] up13_2;
  wire   [4:0] up21_1;
  wire   [4:0] up33_2;
  wire   [4:0] up35_1;
  wire   [4:0] up37_1;
  wire   [4:0] up39_1;
  wire   [4:0] c10_1;
  wire   [4:0] c10_2;
  wire   [4:0] c10_3;
  wire   [4:0] c10_4;
  wire   [4:0] c10_5;
  wire   [4:0] c10_6;
  wire   [4:0] up14_2;
  wire   [4:0] up22_1;
  wire   [4:0] up34_2;
  wire   [4:0] up36_1;
  wire   [4:0] up38_1;
  wire   [4:0] up40_1;
  wire   [4:0] c11_1;
  wire   [4:0] c11_2;
  wire   [4:0] c11_3;
  wire   [4:0] c11_4;
  wire   [4:0] c11_5;
  wire   [4:0] c11_6;
  wire   [4:0] up9_2;
  wire   [4:0] up15_2;
  wire   [4:0] up25_2;
  wire   [4:0] up33_3;
  wire   [4:0] up35_2;
  wire   [4:0] up37_2;
  wire   [4:0] c12_1;
  wire   [4:0] c12_2;
  wire   [4:0] c12_3;
  wire   [4:0] c12_4;
  wire   [4:0] c12_5;
  wire   [4:0] c12_6;
  wire   [4:0] up10_2;
  wire   [4:0] up16_2;
  wire   [4:0] up26_2;
  wire   [4:0] up34_3;
  wire   [4:0] up36_2;
  wire   [4:0] up38_2;
  wire   [4:0] c13_1;
  wire   [4:0] c13_2;
  wire   [4:0] c13_3;
  wire   [4:0] c13_4;
  wire   [4:0] c13_5;
  wire   [4:0] c13_6;
  wire   [4:0] up8_2;
  wire   [4:0] up19_3;
  wire   [4:0] up21_2;
  wire   [4:0] up35_3;
  wire   [4:0] up37_3;
  wire   [4:0] up39_2;
  wire   [4:0] c14_1;
  wire   [4:0] c14_2;
  wire   [4:0] c14_3;
  wire   [4:0] c14_4;
  wire   [4:0] c14_5;
  wire   [4:0] c14_6;
  wire   [4:0] up7_2;
  wire   [4:0] up20_3;
  wire   [4:0] up22_2;
  wire   [4:0] up36_3;
  wire   [4:0] up38_3;
  wire   [4:0] up40_2;
  wire   [4:0] c15_1;
  wire   [4:0] c15_2;
  wire   [4:0] c15_3;
  wire   [4:0] c15_4;
  wire   [4:0] c15_5;
  wire   [4:0] c15_6;
  wire   [4:0] up4_3;
  wire   [4:0] up13_3;
  wire   [4:0] up27_3;
  wire   [4:0] up41_1;
  wire   [4:0] up43_1;
  wire   [4:0] up45_1;
  wire   [4:0] c16_1;
  wire   [4:0] c16_2;
  wire   [4:0] c16_3;
  wire   [4:0] c16_4;
  wire   [4:0] c16_5;
  wire   [4:0] c16_6;
  wire   [4:0] up3_3;
  wire   [4:0] up14_3;
  wire   [4:0] up28_3;
  wire   [4:0] up42_1;
  wire   [4:0] up44_1;
  wire   [4:0] up46_1;
  wire   [4:0] c17_1;
  wire   [4:0] c17_2;
  wire   [4:0] c17_3;
  wire   [4:0] c17_4;
  wire   [4:0] c17_5;
  wire   [4:0] c17_6;
  wire   [4:0] up1_2;
  wire   [4:0] up10_3;
  wire   [4:0] up11_2;
  wire   [4:0] up24_1;
  wire   [4:0] up39_3;
  wire   [4:0] up41_2;
  wire   [4:0] c18_1;
  wire   [4:0] c18_2;
  wire   [4:0] c18_3;
  wire   [4:0] c18_4;
  wire   [4:0] c18_5;
  wire   [4:0] c18_6;
  wire   [4:0] up2_2;
  wire   [4:0] up9_3;
  wire   [4:0] up12_2;
  wire   [4:0] up23_1;
  wire   [4:0] up40_3;
  wire   [4:0] up42_2;
  wire   [4:0] c19_1;
  wire   [4:0] c19_2;
  wire   [4:0] c19_3;
  wire   [4:0] c19_4;
  wire   [4:0] c19_5;
  wire   [4:0] c19_6;
  wire   [4:0] up11_3;
  wire   [4:0] up21_3;
  wire   [4:0] up23_2;
  wire   [4:0] up41_3;
  wire   [4:0] up43_2;
  wire   [4:0] up47_1;
  wire   [4:0] c20_1;
  wire   [4:0] c20_2;
  wire   [4:0] c20_3;
  wire   [4:0] c20_4;
  wire   [4:0] c20_5;
  wire   [4:0] c20_6;
  wire   [4:0] up12_3;
  wire   [4:0] up22_3;
  wire   [4:0] up24_2;
  wire   [4:0] up42_3;
  wire   [4:0] up44_2;
  wire   [4:0] up48_1;
  wire   [4:0] c21_1;
  wire   [4:0] c21_2;
  wire   [4:0] c21_3;
  wire   [4:0] c21_4;
  wire   [4:0] c21_5;
  wire   [4:0] c21_6;
  wire   [4:0] up6_3;
  wire   [4:0] up8_3;
  wire   [4:0] up18_3;
  wire   [4:0] up43_3;
  wire   [4:0] up45_2;
  wire   [4:0] up47_2;
  wire   [4:0] c22_1;
  wire   [4:0] c22_2;
  wire   [4:0] c22_3;
  wire   [4:0] c22_4;
  wire   [4:0] c22_5;
  wire   [4:0] c22_6;
  wire   [4:0] up5_3;
  wire   [4:0] up7_3;
  wire   [4:0] up17_3;
  wire   [4:0] up44_3;
  wire   [4:0] up46_2;
  wire   [4:0] up48_2;
  wire   [4:0] c23_1;
  wire   [4:0] c23_2;
  wire   [4:0] c23_3;
  wire   [4:0] c23_4;
  wire   [4:0] c23_5;
  wire   [4:0] c23_6;
  wire   [4:0] up2_3;
  wire   [4:0] up16_3;
  wire   [4:0] up23_3;
  wire   [4:0] up26_3;
  wire   [4:0] up45_3;
  wire   [4:0] up47_3;
  wire   [4:0] c24_1;
  wire   [4:0] c24_2;
  wire   [4:0] c24_3;
  wire   [4:0] c24_4;
  wire   [4:0] c24_5;
  wire   [4:0] c24_6;
  wire   [4:0] up1_3;
  wire   [4:0] up15_3;
  wire   [4:0] up24_3;
  wire   [4:0] up25_3;
  wire   [4:0] up46_3;

  all6_23 all_1 ( .r1(c1_1), .r2(c1_2), .r3(c1_3), .r4(c1_4), .r5(c1_5), .r6(
        c1_6), .i1(up3_1), .i2(up6_1), .i3({up18_1[4:3], n74, up18_1[1:0]}), 
        .i4(up20_1), .i5(up26_1), .i6(up27_1) );
  all6_22 all_2 ( .r1(c2_1), .r2(c2_2), .r3(c2_3), .r4(c2_4), .r5(c2_5), .r6(
        c2_6), .i1(up4_1), .i2(up5_1), .i3(up17_1), .i4(up19_1), .i5(up25_1), 
        .i6(up28_1) );
  all6_21 all_3 ( .r1(c3_1), .r2(c3_2), .r3(c3_3), .r4(c3_4), .r5(c3_5), .r6(
        c3_6), .i1(up4_2), .i2(up14_1), .i3(up16_1), .i4(up27_2), .i5(up29_1), 
        .i6(up31_1) );
  all6_20 all_4 ( .r1(c4_1), .r2(c4_2), .r3(c4_3), .r4(c4_4), .r5(c4_5), .r6(
        c4_6), .i1(up3_2), .i2(up13_1), .i3(up15_1), .i4(up28_2), .i5(up30_1), 
        .i6(up32_1) );
  all6_19 all_5 ( .r1(c5_1), .r2(c5_2), .r3(c5_3), .r4(c5_4), .r5(c5_5), .r6(
        c5_6), .i1(up7_1), .i2(up9_1), .i3(up12_1), .i4(up29_2), .i5(up31_2), 
        .i6(up33_1) );
  all6_18 all_6 ( .r1(c6_1), .r2(c6_2), .r3(c6_3), .r4(c6_4), .r5(c6_5), .r6(
        c6_6), .i1(up8_1), .i2(up10_1), .i3(up11_1), .i4(up30_2), .i5(up32_2), 
        .i6(up34_1) );
  all6_17 all_7 ( .r1(c7_1), .r2(c7_2), .r3(c7_3), .r4(c7_4), .r5(c7_5), .r6(
        c7_6), .i1(up2_1), .i2(up6_2), .i3(up18_2), .i4(up20_2), .i5(up29_3), 
        .i6(up31_3) );
  all6_16 all_8 ( .r1(c8_1), .r2(c8_2), .r3(c8_3), .r4(c8_4), .r5(c8_5), .r6(
        c8_6), .i1(up1_1), .i2(up5_2), .i3(up17_2), .i4(up19_2), .i5(up30_3), 
        .i6(up32_3) );
  all6_15 all_9 ( .r1(c9_1), .r2(c9_2), .r3(c9_3), .r4(c9_4), .r5(c9_5), .r6(
        c9_6), .i1(up13_2), .i2(up21_1), .i3(up33_2), .i4(up35_1), .i5(up37_1), 
        .i6(up39_1) );
  all6_14 all_10 ( .r1(c10_1), .r2(c10_2), .r3(c10_3), .r4(c10_4), .r5(c10_5), 
        .r6(c10_6), .i1(up14_2), .i2(up22_1), .i3(up34_2), .i4(up36_1), .i5(
        up38_1), .i6(up40_1) );
  all6_13 all_11 ( .r1(c11_1), .r2(c11_2), .r3(c11_3), .r4(c11_4), .r5(c11_5), 
        .r6(c11_6), .i1(up9_2), .i2(up15_2), .i3(up25_2), .i4(up33_3), .i5(
        up35_2), .i6(up37_2) );
  all6_12 all_12 ( .r1(c12_1), .r2(c12_2), .r3(c12_3), .r4(c12_4), .r5(c12_5), 
        .r6(c12_6), .i1(up10_2), .i2(up16_2), .i3(up26_2), .i4({n76, 
        up34_3[3:0]}), .i5(up36_2), .i6(up38_2) );
  all6_11 all_13 ( .r1(c13_1), .r2(c13_2), .r3(c13_3), .r4(c13_4), .r5(c13_5), 
        .r6(c13_6), .i1(up8_2), .i2(up19_3), .i3(up21_2), .i4(up35_3), .i5(
        up37_3), .i6(up39_2) );
  all6_10 all_14 ( .r1(c14_1), .r2(c14_2), .r3(c14_3), .r4(c14_4), .r5(c14_5), 
        .r6(c14_6), .i1(up7_2), .i2(up20_3), .i3(up22_2), .i4(up36_3), .i5(
        up38_3), .i6(up40_2) );
  all6_9 all_15 ( .r1(c15_1), .r2(c15_2), .r3(c15_3), .r4(c15_4), .r5(c15_5), 
        .r6(c15_6), .i1(up4_3), .i2(up13_3), .i3(up27_3), .i4(up41_1), .i5(
        up43_1), .i6(up45_1) );
  all6_8 all_16 ( .r1(c16_1), .r2(c16_2), .r3(c16_3), .r4(c16_4), .r5(c16_5), 
        .r6(c16_6), .i1(up3_3), .i2(up14_3), .i3(up28_3), .i4(up42_1), .i5(
        up44_1), .i6(up46_1) );
  all6_7 all_17 ( .r1(c17_1), .r2(c17_2), .r3(c17_3), .r4(c17_4), .r5(c17_5), 
        .r6(c17_6), .i1(up1_2), .i2(up10_3), .i3({up11_2[4:3], n77, 
        up11_2[1:0]}), .i4(up24_1), .i5(up39_3), .i6(up41_2) );
  all6_6 all_18 ( .r1(c18_1), .r2(c18_2), .r3(c18_3), .r4(c18_4), .r5(c18_5), 
        .r6(c18_6), .i1({n75, up2_2[3:0]}), .i2(up9_3), .i3(up12_2), .i4(
        up23_1), .i5(up40_3), .i6(up42_2) );
  all6_5 all_19 ( .r1(c19_1), .r2(c19_2), .r3(c19_3), .r4(c19_4), .r5(c19_5), 
        .r6(c19_6), .i1({n118, up11_3[3:0]}), .i2(up21_3), .i3(up23_2), .i4(
        up41_3), .i5(up43_2), .i6({up47_1[4:3], n120, up47_1[1:0]}) );
  all6_4 all_20 ( .r1(c20_1), .r2(c20_2), .r3(c20_3), .r4(c20_4), .r5(c20_5), 
        .r6(c20_6), .i1({n117, up12_3[3:0]}), .i2({up22_3[4:1], n78}), .i3(
        up24_2), .i4({n116, up42_3[3:0]}), .i5(up44_2), .i6(up48_1) );
  all6_3 all_21 ( .r1(c21_1), .r2(c21_2), .r3(c21_3), .r4(c21_4), .r5(c21_5), 
        .r6(c21_6), .i1(up6_3), .i2(up8_3), .i3(up18_3), .i4(up43_3), .i5(
        up45_2), .i6(up47_2) );
  all6_2 all_22 ( .r1(c22_1), .r2(c22_2), .r3(c22_3), .r4(c22_4), .r5(c22_5), 
        .r6(c22_6), .i1({n119, up5_3[3:0]}), .i2(up7_3), .i3(up17_3), .i4(
        up44_3), .i5(up46_2), .i6(up48_2) );
  all6_1 all_23 ( .r1(c23_1), .r2(c23_2), .r3(c23_3), .r4(c23_4), .r5(c23_5), 
        .r6(c23_6), .i1(up2_3), .i2(up16_3), .i3(up23_3), .i4(up26_3), .i5(
        up45_3), .i6(up47_3) );
  all6_0 all_24 ( .r1(c24_1), .r2(c24_2), .r3(c24_3), .r4(c24_4), .r5(c24_5), 
        .r6(c24_6), .i1(up1_3), .i2(up15_3), .i3(up24_3), .i4(up25_3), .i5(
        up46_3), .i6({test_so, up48_3_3_, up48_3_2_, up48_3_1_, up48_3_0_}) );
  total_3_test_0 total_1 ( .h(h1), .up1(up1_1), .up2(up1_2), .up3(up1_3), 
        .clk(clk), .rst(n84), .a(c8_1), .b(c17_1), .c(c24_1), .in(i1), 
        .test_si(test_si), .test_se(n88) );
  total_3_test_1 total_2 ( .h(h2), .up1(up2_1), .up2(up2_2), .up3(up2_3), 
        .clk(clk), .rst(n84), .a({c7_1[4:2], n87, c7_1[0]}), .b(c18_1), .c(
        c23_1), .in(i2), .test_si(up1_3[4]), .test_se(n89) );
  total_3_test_2 total_3 ( .h(h3), .up1(up3_1), .up2(up3_2), .up3(up3_3), 
        .clk(clk), .rst(n84), .a(c1_1), .b(c4_1), .c(c16_1), .in(i3), 
        .test_si(up2_3[4]), .test_se(n90) );
  total_3_test_3 total_4 ( .h(h4), .up1(up4_1), .up2(up4_2), .up3(up4_3), 
        .clk(clk), .rst(n84), .a(c2_1), .b(c3_1), .c(c15_1), .in(i4), 
        .test_si(up3_3[4]), .test_se(n91) );
  total_3_test_4 total_5 ( .h(h5), .up1(up5_1), .up2(up5_2), .up3(up5_3), 
        .clk(clk), .rst(n84), .a(c2_2), .b(c8_2), .c(c22_1), .in(i5), 
        .test_si(up4_3[4]), .test_se(n88) );
  total_3_test_5 total_6 ( .h(h6), .up1(up6_1), .up2(up6_2), .up3(up6_3), 
        .clk(clk), .rst(n84), .a(c1_2), .b(c7_2), .c(c21_1), .in(i6), 
        .test_si(n119), .test_se(n89) );
  total_3_test_6 total_7 ( .h(h7), .up1(up7_1), .up2(up7_2), .up3(up7_3), 
        .clk(clk), .rst(n84), .a(c5_1), .b(c14_1), .c(c22_2), .in(i7), 
        .test_si(up6_3[4]), .test_se(n90) );
  total_3_test_7 total_8 ( .h(h8), .up1(up8_1), .up2(up8_2), .up3(up8_3), 
        .clk(clk), .rst(n84), .a(c6_1), .b(c13_1), .c(c21_2), .in(i8), 
        .test_si(up7_3[4]), .test_se(n91) );
  total_3_test_8 total_9 ( .h(h9), .up1(up9_1), .up2(up9_2), .up3(up9_3), 
        .clk(clk), .rst(n84), .a(c5_2), .b(c11_1), .c(c18_2), .in(i9), 
        .test_si(up8_3[4]), .test_se(n92) );
  total_3_test_9 total_10 ( .h(h10), .up1(up10_1), .up2(up10_2), .up3(up10_3), 
        .clk(clk), .rst(n84), .a(c6_2), .b(c12_1), .c({c17_2[4], n73, 
        c17_2[2:0]}), .in(i10), .test_si(up9_3[4]), .test_se(n92) );
  total_3_test_10 total_11 ( .h(h11), .up1(up11_1), .up2(up11_2), .up3(up11_3), 
        .clk(clk), .rst(n84), .a(c6_3), .b(c17_3), .c(c19_1), .in(i11), 
        .test_si(up10_3[4]), .test_se(n93) );
  total_3_test_11 total_12 ( .h(h12), .up1(up12_1), .up2(up12_2), .up3(up12_3), 
        .clk(clk), .rst(n84), .a(c5_3), .b(c18_3), .c(c20_1), .in(i12), 
        .test_si(n118), .test_se(n93) );
  total_3_test_12 total_13 ( .h(h13), .up1(up13_1), .up2(up13_2), .up3(up13_3), 
        .clk(clk), .rst(n83), .a(c4_2), .b(c9_1), .c(c15_2), .in(i13), 
        .test_si(n117), .test_se(n94) );
  total_3_test_13 total_14 ( .h(h14), .up1(up14_1), .up2(up14_2), .up3(up14_3), 
        .clk(clk), .rst(n83), .a(c3_2), .b(c10_1), .c(c16_2), .in(i14), 
        .test_si(up13_3[4]), .test_se(n94) );
  total_3_test_14 total_15 ( .h(h15), .up1(up15_1), .up2(up15_2), .up3(up15_3), 
        .clk(clk), .rst(n83), .a(c4_3), .b(c11_2), .c(c24_2), .in(i15), 
        .test_si(up14_3[4]), .test_se(n95) );
  total_3_test_15 total_16 ( .h(h16), .up1(up16_1), .up2(up16_2), .up3(up16_3), 
        .clk(clk), .rst(n83), .a(c3_3), .b(c12_2), .c(c23_2), .in(i16), 
        .test_si(up15_3[4]), .test_se(n95) );
  total_3_test_16 total_17 ( .h(h17), .up1(up17_1), .up2(up17_2), .up3(up17_3), 
        .clk(clk), .rst(n83), .a(c2_3), .b(c8_3), .c(c22_3), .in(i17), 
        .test_si(up16_3[4]), .test_se(n114) );
  total_3_test_17 total_18 ( .h(h18), .up1(up18_1), .up2(up18_2), .up3(up18_3), 
        .clk(clk), .rst(n83), .a(c1_3), .b(c7_3), .c(c21_3), .in(i18), 
        .test_si(up17_3[4]), .test_se(n111) );
  total_3_test_18 total_19 ( .h(h19), .up1(up19_1), .up2(up19_2), .up3(up19_3), 
        .clk(clk), .rst(n83), .a(c2_4), .b({n69, n72, c8_4[2:0]}), .c(c13_2), 
        .in(i19), .test_si(up18_3[4]), .test_se(n101) );
  total_3_test_19 total_20 ( .h(h20), .up1(up20_1), .up2(up20_2), .up3(up20_3), 
        .clk(clk), .rst(n83), .a(c1_4), .b(c7_4), .c(c14_2), .in(i20), 
        .test_si(up19_3[4]), .test_se(n111) );
  total_3_test_20 total_21 ( .h(h21), .up1(up21_1), .up2(up21_2), .up3(up21_3), 
        .clk(clk), .rst(n83), .a(c9_2), .b(c13_3), .c(c19_2), .in(i21), 
        .test_si(up20_3[4]), .test_se(n113) );
  total_3_test_21 total_22 ( .h(h22), .up1(up22_1), .up2(up22_2), .up3(up22_3), 
        .clk(clk), .rst(n83), .a(c10_2), .b(c14_3), .c(c20_2), .in(i22), 
        .test_si(up21_3[4]), .test_se(n111) );
  total_3_test_22 total_23 ( .h(h23), .up1(up23_1), .up2(up23_2), .up3(up23_3), 
        .clk(clk), .rst(n83), .a(c18_4), .b(c19_3), .c(c23_3), .in(i23), 
        .test_si(up22_3[4]), .test_se(n113) );
  total_3_test_23 total_24 ( .h(h24), .up1(up24_1), .up2(up24_2), .up3(up24_3), 
        .clk(clk), .rst(n83), .a(c17_4), .b(c20_3), .c(c24_3), .in(i24), 
        .test_si(up23_3[4]), .test_se(n101) );
  total_3_test_24 total_25 ( .h(h25), .up1(up25_1), .up2(up25_2), .up3(up25_3), 
        .clk(clk), .rst(n82), .a(c2_5), .b(c11_3), .c(c24_4), .in(i25), 
        .test_si(up24_3[4]), .test_se(n113) );
  total_3_test_25 total_26 ( .h(h26), .up1(up26_1), .up2(up26_2), .up3(up26_3), 
        .clk(clk), .rst(n82), .a(c1_5), .b(c12_3), .c(c23_4), .in(i26), 
        .test_si(up25_3[4]), .test_se(n114) );
  total_3_test_26 total_27 ( .h(h27), .up1(up27_1), .up2(up27_2), .up3(up27_3), 
        .clk(clk), .rst(n82), .a(c1_6), .b(c3_4), .c(c15_3), .in(i27), 
        .test_si(up26_3[4]), .test_se(n110) );
  total_3_test_27 total_28 ( .h(h28), .up1(up28_1), .up2(up28_2), .up3(up28_3), 
        .clk(clk), .rst(n82), .a(c2_6), .b(c4_4), .c(c16_3), .in(i28), 
        .test_si(up27_3[4]), .test_se(n98) );
  total_3_test_28 total_29 ( .h(h29), .up1(up29_1), .up2(up29_2), .up3(up29_3), 
        .clk(clk), .rst(n82), .a(c3_5), .b(c5_4), .c(c7_5), .in(i29), 
        .test_si(up28_3[4]), .test_se(n103) );
  total_3_test_29 total_30 ( .h(h30), .up1(up30_1), .up2(up30_2), .up3(up30_3), 
        .clk(clk), .rst(n82), .a(c4_5), .b(c6_4), .c(c8_5), .in(i30), 
        .test_si(up29_3[4]), .test_se(n104) );
  total_3_test_30 total_31 ( .h(h31), .up1(up31_1), .up2(up31_2), .up3(up31_3), 
        .clk(clk), .rst(n82), .a(c3_6), .b(c5_5), .c(c7_6), .in(i31), 
        .test_si(up30_3[4]), .test_se(n105) );
  total_3_test_31 total_32 ( .h(h32), .up1(up32_1), .up2(up32_2), .up3(up32_3), 
        .clk(clk), .rst(n82), .a(c4_6), .b(c6_5), .c(c8_6), .in(i32), 
        .test_si(up31_3[4]), .test_se(n102) );
  total_3_test_32 total_33 ( .h(h33), .up1(up33_1), .up2(up33_2), .up3(up33_3), 
        .clk(clk), .rst(n82), .a(c5_6), .b(c9_3), .c(c11_4), .in(i33), 
        .test_si(up32_3[4]), .test_se(n99) );
  total_3_test_33 total_34 ( .h(h34), .up1(up34_1), .up2(up34_2), .up3(up34_3), 
        .clk(clk), .rst(n82), .a(c6_6), .b(c10_3), .c(c12_4), .in(i34), 
        .test_si(up33_3[4]), .test_se(n99) );
  total_3_test_34 total_35 ( .h(h35), .up1(up35_1), .up2(up35_2), .up3(up35_3), 
        .clk(clk), .rst(n82), .a(c9_4), .b(c11_5), .c(c13_4), .in(i35), 
        .test_si(up34_3[4]), .test_se(n106) );
  total_3_test_35 total_36 ( .h(h36), .up1(up36_1), .up2(up36_2), .up3(up36_3), 
        .clk(clk), .rst(n82), .a(c10_4), .b(c12_5), .c(c14_4), .in(i36), 
        .test_si(up35_3[4]), .test_se(n107) );
  total_3_test_36 total_37 ( .h(h37), .up1(up37_1), .up2(up37_2), .up3(up37_3), 
        .clk(clk), .rst(n80), .a(c9_5), .b({c11_6[4:1], n79}), .c(c13_5), .in(
        i37), .test_si(up36_3[4]), .test_se(n108) );
  total_3_test_37 total_38 ( .h(h38), .up1(up38_1), .up2(up38_2), .up3(up38_3), 
        .clk(clk), .rst(n84), .a(c10_5), .b(c12_6), .c(c14_5), .in(i38), 
        .test_si(up37_3[4]), .test_se(n108) );
  total_3_test_38 total_39 ( .h(h39), .up1(up39_1), .up2(up39_2), .up3(up39_3), 
        .clk(clk), .rst(n81), .a(c9_6), .b({n70, c13_6[3:0]}), .c(c17_5), .in(
        i39), .test_si(up38_3[4]), .test_se(n109) );
  total_3_test_39 total_40 ( .h(h40), .up1(up40_1), .up2(up40_2), .up3(up40_3), 
        .clk(clk), .rst(n83), .a(c10_6), .b(c14_6), .c(c18_5), .in(i40), 
        .test_si(up39_3[4]), .test_se(n110) );
  total_3_test_40 total_41 ( .h(h41), .up1(up41_1), .up2(up41_2), .up3(up41_3), 
        .clk(clk), .rst(n82), .a(c15_4), .b(c17_6), .c(c19_4), .in(i41), 
        .test_si(up40_3[4]), .test_se(n110) );
  total_3_test_41 total_42 ( .h(h42), .up1(up42_1), .up2(up42_2), .up3(up42_3), 
        .clk(clk), .rst(n84), .a(c16_4), .b(c18_6), .c(c20_4), .in(i42), 
        .test_si(up41_3[4]), .test_se(n107) );
  total_3_test_42 total_43 ( .h(h43), .up1(up43_1), .up2(up43_2), .up3(up43_3), 
        .clk(clk), .rst(n83), .a(c15_5), .b(c19_5), .c(c21_4), .in(i43), 
        .test_si(n116), .test_se(n96) );
  total_3_test_43 total_44 ( .h(h44), .up1(up44_1), .up2(up44_2), .up3(up44_3), 
        .clk(clk), .rst(n82), .a(c16_5), .b(c20_5), .c(c22_4), .in(i44), 
        .test_si(up43_3[4]), .test_se(n108) );
  total_3_test_44 total_45 ( .h(h45), .up1(up45_1), .up2(up45_2), .up3(up45_3), 
        .clk(clk), .rst(n84), .a(c15_6), .b(c21_5), .c(c23_5), .in(i45), 
        .test_si(up44_3[4]), .test_se(n97) );
  total_3_test_45 total_46 ( .h(h46), .up1(up46_1), .up2(up46_2), .up3(up46_3), 
        .clk(clk), .rst(n83), .a(c16_6), .b(c22_5), .c(c24_5), .in(i46), 
        .test_si(up45_3[4]), .test_se(n106) );
  total_3_test_46 total_47 ( .h(h47), .up1(up47_1), .up2(up47_2), .up3(up47_3), 
        .clk(clk), .rst(n82), .a(c19_6), .b(c21_6), .c(c23_6), .in(i47), 
        .test_si(up46_3[4]), .test_se(n106) );
  total_3_test_47 total_48 ( .h(h48), .up1(up48_1), .up2(up48_2), .up3({
        test_so, up48_3_3_, up48_3_2_, up48_3_1_, up48_3_0_}), .clk(clk), 
        .rst(n84), .a(c20_6), .b(c22_6), .c(c24_6), .in(i48), .test_si(
        up47_3[4]), .test_se(n107) );
  BUFX2 U1 ( .A(c8_4[4]), .Y(n69) );
  BUFX6 U2 ( .A(up34_3[4]), .Y(n76) );
  CLKBUFX2TH U3 ( .A(c13_6[4]), .Y(n70) );
  BUFX2TH U4 ( .A(up2_2[4]), .Y(n75) );
  BUFX3TH U5 ( .A(c11_6[0]), .Y(n79) );
  INVXLTH U6 ( .A(c8_4[3]), .Y(n71) );
  INVXLTH U7 ( .A(n71), .Y(n72) );
  CLKBUFX1TH U8 ( .A(c17_2[3]), .Y(n73) );
  CLKBUFX2TH U9 ( .A(up18_1[2]), .Y(n74) );
  CLKBUFX2TH U10 ( .A(up11_2[2]), .Y(n77) );
  CLKBUFX2TH U11 ( .A(up22_3[0]), .Y(n78) );
  CLKBUFX1TH U12 ( .A(rst), .Y(n80) );
  CLKBUFX1TH U13 ( .A(rst), .Y(n81) );
  CLKBUFX8TH U14 ( .A(n80), .Y(n82) );
  CLKBUFX8TH U15 ( .A(n81), .Y(n83) );
  CLKBUFX8TH U16 ( .A(n81), .Y(n84) );
  CLKBUFX40 U17 ( .A(c7_1[1]), .Y(n87) );
  DLY1X1TH U18 ( .A(test_se), .Y(n88) );
  DLY1X1TH U19 ( .A(test_se), .Y(n89) );
  DLY1X1TH U20 ( .A(test_se), .Y(n90) );
  DLY1X1TH U21 ( .A(test_se), .Y(n91) );
  DLY1X1TH U22 ( .A(n88), .Y(n92) );
  DLY1X1TH U23 ( .A(n92), .Y(n93) );
  DLY1X1TH U24 ( .A(n93), .Y(n94) );
  DLY1X1TH U25 ( .A(n94), .Y(n95) );
  DLY1X1TH U26 ( .A(n97), .Y(n96) );
  DLY1X1TH U27 ( .A(n98), .Y(n97) );
  DLY1X1TH U28 ( .A(n102), .Y(n98) );
  DLY1X1TH U29 ( .A(n104), .Y(n99) );
  DLY1X1TH U30 ( .A(n112), .Y(n100) );
  DLY1X1TH U31 ( .A(n112), .Y(n101) );
  DLY1X1TH U32 ( .A(n115), .Y(n102) );
  DLY1X1TH U33 ( .A(n115), .Y(n103) );
  DLY1X1TH U34 ( .A(n115), .Y(n104) );
  DLY1X1TH U35 ( .A(n115), .Y(n105) );
  DLY1X1TH U36 ( .A(n98), .Y(n106) );
  DLY1X1TH U37 ( .A(n103), .Y(n107) );
  DLY1X1TH U38 ( .A(n114), .Y(n108) );
  DLY1X1TH U39 ( .A(n100), .Y(n109) );
  DLY1X1TH U40 ( .A(n112), .Y(n110) );
  DLY1X1TH U41 ( .A(n112), .Y(n111) );
  DLY1X1TH U42 ( .A(n95), .Y(n112) );
  DLY1X1TH U43 ( .A(n100), .Y(n113) );
  DLY1X1TH U44 ( .A(n100), .Y(n114) );
  DLY1X1TH U45 ( .A(n101), .Y(n115) );
  DLY1X1TH U46 ( .A(up42_3[4]), .Y(n116) );
  DLY1X1TH U47 ( .A(up12_3[4]), .Y(n117) );
  DLY1X1TH U48 ( .A(up11_3[4]), .Y(n118) );
  DLY1X1TH U49 ( .A(up5_3[4]), .Y(n119) );
  CLKBUFX40 U50 ( .A(up47_1[2]), .Y(n120) );
endmodule


module data_mux ( out, in1, in2, sel );
  output [4:0] out;
  input [4:0] in1;
  input [4:0] in2;
  input sel;
  wire   n2;

  CLKINVX2TH U1 ( .A(sel), .Y(n2) );
  AO22XLTH U2 ( .A0(in2[4]), .A1(n2), .B0(sel), .B1(in1[4]), .Y(out[4]) );
  AO22XLTH U3 ( .A0(in2[1]), .A1(n2), .B0(in1[1]), .B1(sel), .Y(out[1]) );
  AO22XLTH U4 ( .A0(in2[3]), .A1(n2), .B0(in1[3]), .B1(sel), .Y(out[3]) );
  AO22XLTH U5 ( .A0(in2[0]), .A1(n2), .B0(in1[0]), .B1(sel), .Y(out[0]) );
  AO22XLTH U6 ( .A0(in2[2]), .A1(n2), .B0(in1[2]), .B1(sel), .Y(out[2]) );
endmodule


module segma_table ( out, in );
  output [15:0] out;
  input [2:0] in;
  wire   n6, n7, n8, n24, n25, n26, n27;

  INVX2TH U3 ( .A(1'b0), .Y(out[14]) );
  INVX2TH U5 ( .A(1'b1), .Y(out[15]) );
  AOI2BB1XLTH U7 ( .A0N(in[1]), .A1N(n27), .B0(in[2]), .Y(out[2]) );
  NAND2X1TH U8 ( .A(in[2]), .B(in[1]), .Y(out[13]) );
  OAI221XLTH U9 ( .A0(in[0]), .A1(out[13]), .B0(in[2]), .B1(n27), .C0(n25), 
        .Y(out[11]) );
  NOR2X1TH U10 ( .A(in[1]), .B(in[2]), .Y(out[6]) );
  OAI211XLTH U11 ( .A0(in[0]), .A1(n24), .B0(n8), .C0(n25), .Y(out[7]) );
  NAND2XLTH U12 ( .A(in[1]), .B(in[0]), .Y(n8) );
  CLKINVX1TH U13 ( .A(in[2]), .Y(n24) );
  CLKXOR2X2TH U14 ( .A(in[1]), .B(in[0]), .Y(n6) );
  INVXLTH U15 ( .A(out[6]), .Y(n25) );
  CLKINVX1TH U16 ( .A(in[0]), .Y(n27) );
  CLKINVX1TH U17 ( .A(n8), .Y(n26) );
  NAND2BX1TH U18 ( .AN(n6), .B(n24), .Y(n7) );
  OAI21XLTH U19 ( .A0(in[2]), .A1(n26), .B0(out[13]), .Y(out[12]) );
  CLKBUFX1TH U20 ( .A(out[6]), .Y(out[3]) );
  NOR2XLTH U21 ( .A(n26), .B(n7), .Y(out[0]) );
  OAI21XLTH U22 ( .A0(in[0]), .A1(out[13]), .B0(n7), .Y(out[1]) );
  AOI21XLTH U23 ( .A0(n26), .A1(n24), .B0(n6), .Y(out[10]) );
  INVXLTH U26 ( .A(n6), .Y(out[8]) );
  OAI21XLTH U27 ( .A0(n26), .A1(n6), .B0(n7), .Y(out[5]) );
  NAND2XLTH U28 ( .A(in[2]), .B(n6), .Y(out[4]) );
  AO21XLTH U29 ( .A0(n27), .A1(in[1]), .B0(out[2]), .Y(out[9]) );
endmodule


module multiplier_1_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;
  wire   n2, n3;
  wire   [15:3] carry;

  XOR2X1 U1 ( .A(A[11]), .B(carry[11]), .Y(SUM[11]) );
  ADDHX2 U1_1_12 ( .A(A[12]), .B(n3), .CO(carry[13]), .S(SUM[12]) );
  ADDHX1TH U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXLTH U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHX4 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHX2 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHX1TH U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHX1 U1_1_2 ( .A(A[2]), .B(n2), .CO(carry[3]), .S(SUM[2]) );
  ADDHX1TH U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX2 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHX4 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  CLKAND2X4 U2 ( .A(A[11]), .B(carry[11]), .Y(n3) );
  XOR2X1 U3 ( .A(A[1]), .B(A[0]), .Y(SUM[1]) );
  AND2XLTH U4 ( .A(A[1]), .B(A[0]), .Y(n2) );
  INVXLTH U5 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X8 U6 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
endmodule


module multiplier_1_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  ADDHX1TH U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHX2TH U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHX4 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHX4 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHX4 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHX4 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4TH U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHX4TH U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4TH U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHX2 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHX2 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHX2TH U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  INVX2TH U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module multiplier_1_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;
  wire   n1, n5, n6, n7, n8;
  wire   [15:2] carry;

  ADDHX4 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHX4 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHX4 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX2TH U1_1_5 ( .A(A[5]), .B(n1), .CO(carry[6]), .S(SUM[5]) );
  ADDHX2TH U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHX2 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHX2 U1_1_12 ( .A(A[12]), .B(n7), .CO(carry[13]), .S(SUM[12]) );
  ADDHX2 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHX4 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHX2 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  XOR2X4 U1 ( .A(A[11]), .B(carry[11]), .Y(SUM[11]) );
  CLKAND2X4 U2 ( .A(A[4]), .B(carry[4]), .Y(n1) );
  AND2XLTH U3 ( .A(A[11]), .B(carry[11]), .Y(n7) );
  XOR2X1 U4 ( .A(A[4]), .B(carry[4]), .Y(SUM[4]) );
  CLKNAND2X2 U5 ( .A(n5), .B(n6), .Y(SUM[15]) );
  NAND2BX2TH U6 ( .AN(carry[15]), .B(A[15]), .Y(n6) );
  NAND2XLTH U7 ( .A(carry[15]), .B(n8), .Y(n5) );
  INVXLTH U8 ( .A(A[0]), .Y(SUM[0]) );
  INVXLTH U9 ( .A(A[15]), .Y(n8) );
endmodule


module multiplier_1_DW_mult_uns_3 ( a, b, product_30_, product_29_, 
        product_28_, product_27_, product_26_, product_25_, product_24_, 
        product_23_, product_22_, product_21_, product_20_, product_19_, 
        product_18_, product_17_, product_16_, product_15_ );
  input [15:0] a;
  input [15:0] b;
  output product_30_, product_29_, product_28_, product_27_, product_26_,
         product_25_, product_24_, product_23_, product_22_, product_21_,
         product_20_, product_19_, product_18_, product_17_, product_16_,
         product_15_;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n68, n70, n71, n72, n76, n77, n78, n79, n80, n84, n85, n86,
         n87, n88, n92, n93, n94, n95, n96, n100, n101, n102, n103, n104, n108,
         n109, n110, n111, n112, n116, n117, n118, n119, n120, n124, n125,
         n126, n127, n128, n132, n134, n135, n136, n139, n140, n147, n148,
         n155, n156, n158, n159, n160, n163, n166, n171, n172, n174, n175,
         n176, n179, n182, n199, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n773, n774, n775, n777, n778,
         n779, n780, n781, n784, n785, n787, n791, n793, n795, n796, n864,
         n865, n866, n867, n868, n871, n872, n874, n875, n876, n877, n880,
         n881, n882, n883, n884, n885, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n906, n907, n908, n909, n910, n911, n912, n914, n915, n916,
         n917, n918, n919, n925, n926, n927, n928, n929, n930, n932, n933,
         n936, n937, n938, n939, n940, n946, n947, n949, n950, n951, n954,
         n955, n957, n958, n959, n960, n961, n962, n964, n965, n966, n967,
         n969, n970, n977, n978, n983, n987, n988, n989, n990, n991, n992,
         n993, n994, n1019, n1020, n1021, n1022, n1024, n1027, n1028, n1029,
         n1030, n1031, n1034, n1035, n1038, n1039, n1041, n1042, n1049, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191;

  OAI22X1 U1095 ( .A0(n1147), .A1(n735), .B0(n734), .B1(n796), .Y(n586) );
  XNOR2X1 U850 ( .A(n1143), .B(n1074), .Y(n659) );
  NAND2X2 U994 ( .A(n957), .B(n958), .Y(n774) );
  XNOR2X1 U1058 ( .A(n1142), .B(n1061), .Y(n687) );
  OAI22X1 U1405 ( .A0(n785), .A1(n704), .B0(n703), .B1(n1096), .Y(n553) );
  OAI22X1 U779 ( .A0(n1146), .A1(n1089), .B0(n688), .B1(n793), .Y(n451) );
  NAND2X2 U1128 ( .A(n292), .B(n305), .Y(n111) );
  NAND2X2 U1272 ( .A(n1144), .B(n1168), .Y(n957) );
  NAND2X2 U1281 ( .A(n914), .B(n915), .Y(n684) );
  NAND2BX2 U1336 ( .AN(n1061), .B(n1143), .Y(n671) );
  NAND2BX2 U1478 ( .AN(n1061), .B(n1142), .Y(n688) );
  NAND3X2 U707 ( .A(n917), .B(n918), .C(n919), .Y(n293) );
  ADDFX1 U708 ( .A(n313), .B(n300), .CI(n298), .CO(n295), .S(n296) );
  CLKXOR2X4 U709 ( .A(n889), .B(n302), .Y(n300) );
  CLKNAND2X4 U710 ( .A(n946), .B(n947), .Y(n775) );
  XNOR2X1 U711 ( .A(n109), .B(n61), .Y(product_20_) );
  NAND2X4 U712 ( .A(n1112), .B(n111), .Y(n109) );
  CLKNAND2X8 U713 ( .A(n85), .B(n926), .Y(n1110) );
  OAI21X6 U714 ( .A0(n88), .A1(n86), .B0(n87), .Y(n85) );
  OAI21X4 U715 ( .A0(n120), .A1(n118), .B0(n119), .Y(n117) );
  CLKNAND2X2 U716 ( .A(n322), .B(n336), .Y(n119) );
  AOI21BX2 U717 ( .A0(n125), .A1(n1049), .B0N(n124), .Y(n120) );
  AND2X2 U718 ( .A(n951), .B(n132), .Y(n128) );
  NAND2BX8 U719 ( .AN(n993), .B(n1098), .Y(n951) );
  CLKXOR2X2 U720 ( .A(n565), .B(n549), .Y(n407) );
  XOR3X2 U721 ( .A(n388), .B(n381), .C(n390), .Y(n377) );
  ADDFX4 U722 ( .A(n393), .B(n400), .CI(n391), .CO(n388), .S(n389) );
  ADDFHX2 U723 ( .A(n599), .B(n536), .CI(n552), .CO(n426), .S(n427) );
  OAI22XL U724 ( .A0(n785), .A1(n703), .B0(n702), .B1(n1096), .Y(n552) );
  OR2X8 U725 ( .A(n365), .B(n376), .Y(n1098) );
  ADDFHX4 U726 ( .A(n369), .B(n378), .CI(n367), .CO(n364), .S(n365) );
  BUFX6 U727 ( .A(a[4]), .Y(n1054) );
  CLKNAND2X2 U728 ( .A(a[8]), .B(n1141), .Y(n1024) );
  XNOR2X4 U729 ( .A(n1142), .B(a[8]), .Y(n1101) );
  BUFX6 U730 ( .A(n749), .Y(n1055) );
  XNOR2XL U731 ( .A(n1130), .B(n1138), .Y(n749) );
  NAND2BX2 U732 ( .AN(n1152), .B(n124), .Y(n65) );
  CLKNAND2X2 U733 ( .A(n337), .B(n350), .Y(n124) );
  INVX4 U734 ( .A(a[8]), .Y(n1174) );
  OAI22XL U735 ( .A0(n785), .A1(n702), .B0(n701), .B1(n1095), .Y(n551) );
  XNOR2XL U736 ( .A(n1137), .B(n1140), .Y(n706) );
  BUFX12 U737 ( .A(b[15]), .Y(n1137) );
  OAI22X2 U738 ( .A0(n744), .A1(n1125), .B0(n745), .B1(n1069), .Y(n596) );
  OAI22X2 U739 ( .A0(n743), .A1(n1125), .B0(n744), .B1(n1069), .Y(n595) );
  XNOR2X1 U740 ( .A(n1074), .B(n1138), .Y(n744) );
  BUFX20 U741 ( .A(b[1]), .Y(n1056) );
  ADDFHX2 U742 ( .A(n501), .B(n380), .CI(n371), .CO(n366), .S(n367) );
  OAI22XL U743 ( .A0(n1077), .A1(n652), .B0(n651), .B1(n791), .Y(n501) );
  ADDFHX2 U744 ( .A(n360), .B(n576), .CI(n499), .CO(n344), .S(n345) );
  OAI22XL U745 ( .A0(n1077), .A1(n650), .B0(n649), .B1(n791), .Y(n499) );
  ADDFHX1 U746 ( .A(n348), .B(n498), .CI(n346), .CO(n329), .S(n330) );
  CLKBUFX40 U747 ( .A(a[3]), .Y(n1139) );
  BUFX3 U748 ( .A(n1164), .Y(n1057) );
  BUFX5 U749 ( .A(n1164), .Y(n1058) );
  BUFX16 U750 ( .A(n1164), .Y(n1059) );
  INVX2 U751 ( .A(n1145), .Y(n1164) );
  ADDFHX1 U752 ( .A(n502), .B(n449), .CI(n383), .CO(n378), .S(n379) );
  OAI22X2 U753 ( .A0(n1062), .A1(n716), .B0(n715), .B1(n795), .Y(n566) );
  OAI22X4 U754 ( .A0(n714), .A1(n795), .B0(n1062), .B1(n715), .Y(n565) );
  XNOR2X1 U755 ( .A(n1130), .B(n1140), .Y(n715) );
  NAND2X6 U756 ( .A(n1093), .B(n1094), .Y(n743) );
  ADDFHX2 U757 ( .A(n558), .B(n497), .CI(n331), .CO(n313), .S(n314) );
  OAI22XL U758 ( .A0(n1077), .A1(n648), .B0(n647), .B1(n791), .Y(n497) );
  NAND2XL U759 ( .A(n496), .B(n317), .Y(n892) );
  XOR2X4 U760 ( .A(n317), .B(n496), .Y(n889) );
  CLKNAND2X2 U761 ( .A(n302), .B(n496), .Y(n890) );
  OAI22X1 U762 ( .A0(n1077), .A1(n647), .B0(n646), .B1(n791), .Y(n496) );
  OAI22X2 U763 ( .A0(n732), .A1(n796), .B0(n733), .B1(n1147), .Y(n584) );
  XNOR2X1 U764 ( .A(n1130), .B(n1139), .Y(n732) );
  BUFX16 U765 ( .A(b[10]), .Y(n1134) );
  NOR2BX8 U766 ( .AN(n1148), .B(n1103), .Y(n519) );
  OAI22X2TH U767 ( .A0(n1073), .A1(n664), .B0(n663), .B1(n1103), .Y(n512) );
  OAI22X4 U768 ( .A0(n1073), .A1(n669), .B0(n668), .B1(n1103), .Y(n517) );
  OAI22X1 U769 ( .A0(n1073), .A1(n670), .B0(n669), .B1(n1103), .Y(n518) );
  CLKNAND2X12 U770 ( .A(n1090), .B(n1091), .Y(n1103) );
  ADDFHX2 U771 ( .A(n580), .B(n532), .CI(n397), .CO(n394), .S(n395) );
  OAI22X1 U772 ( .A0(n728), .A1(n796), .B0(n729), .B1(n1147), .Y(n580) );
  XNOR2X4 U773 ( .A(n1138), .B(n1126), .Y(n753) );
  XNOR2X4 U774 ( .A(n1140), .B(n1126), .Y(n719) );
  XNOR2X4 U775 ( .A(n1139), .B(n1126), .Y(n736) );
  XNOR2X4 U776 ( .A(n1141), .B(n1126), .Y(n702) );
  XNOR2X4 U777 ( .A(n1142), .B(n1126), .Y(n685) );
  XNOR2X1 U778 ( .A(n1143), .B(n1126), .Y(n668) );
  BUFX12 U780 ( .A(b[2]), .Y(n1126) );
  BUFX14 U781 ( .A(b[0]), .Y(n1060) );
  CLKBUFX12 U782 ( .A(b[0]), .Y(n1061) );
  CLKBUFX40 U783 ( .A(a[7]), .Y(n1141) );
  INVX2 U784 ( .A(n1135), .Y(n1182) );
  BUFX20 U785 ( .A(b[13]), .Y(n1135) );
  BUFX20 U786 ( .A(n1076), .Y(n1062) );
  NAND2X8 U787 ( .A(n778), .B(n795), .Y(n1076) );
  INVX20 U788 ( .A(n1131), .Y(n1186) );
  BUFX20 U789 ( .A(b[7]), .Y(n1131) );
  ADDFX2 U790 ( .A(n564), .B(n548), .CI(n929), .CO(n396), .S(n397) );
  NAND2X5 U791 ( .A(n1041), .B(n1042), .Y(n714) );
  BUFX10 U792 ( .A(n585), .Y(n1063) );
  BUFX4 U793 ( .A(a[2]), .Y(n1064) );
  BUFX5 U794 ( .A(n454), .Y(n1065) );
  NAND2XL U795 ( .A(n1138), .B(n1125), .Y(n969) );
  NAND2X4 U796 ( .A(n780), .B(n1125), .Y(n1075) );
  OAI22X4 U797 ( .A0(n1069), .A1(n755), .B0(n754), .B1(n1125), .Y(n606) );
  OAI22X4 U798 ( .A0(n1069), .A1(n1179), .B0(n756), .B1(n1125), .Y(n455) );
  CLKBUFX40 U799 ( .A(n1158), .Y(n1125) );
  OAI22XL U800 ( .A0(n693), .A1(n1096), .B0(n694), .B1(n785), .Y(n543) );
  NAND2X1 U801 ( .A(n1179), .B(a[0]), .Y(n970) );
  OAI22XL U802 ( .A0(n711), .A1(n795), .B0(n712), .B1(n1062), .Y(n562) );
  OAI22XL U803 ( .A0(n781), .A1(n1059), .B0(n637), .B1(n1066), .Y(n448) );
  OAI22X1 U804 ( .A0(n781), .A1(n636), .B0(n635), .B1(n1066), .Y(n485) );
  ADDFX2 U805 ( .A(n387), .B(n531), .CI(n579), .CO(n384), .S(n385) );
  ADDFHX2 U806 ( .A(n514), .B(n577), .CI(n361), .CO(n358), .S(n359) );
  NOR2X1 U807 ( .A(n1058), .B(n1189), .Y(n466) );
  OAI22XL U808 ( .A0(n781), .A1(n634), .B0(n633), .B1(n1066), .Y(n483) );
  INVX2TH U809 ( .A(n126), .Y(n1153) );
  OAI22XLTH U810 ( .A0(n1147), .A1(n1177), .B0(n739), .B1(n796), .Y(n454) );
  CLKNAND2X2 U811 ( .A(n880), .B(n881), .Y(n735) );
  OAI22X1 U812 ( .A0(n733), .A1(n796), .B0(n1147), .B1(n734), .Y(n585) );
  NAND2XLTH U813 ( .A(n571), .B(n443), .Y(n960) );
  NOR2X2TH U814 ( .A(n1099), .B(n166), .Y(n897) );
  NOR2X2TH U815 ( .A(n785), .B(n698), .Y(n898) );
  XNOR2X1TH U816 ( .A(n1072), .B(n1139), .Y(n726) );
  XNOR2X1TH U817 ( .A(n1072), .B(n1142), .Y(n675) );
  BUFX8 U818 ( .A(b[6]), .Y(n1130) );
  BUFX5 U819 ( .A(b[8]), .Y(n1132) );
  CLKNAND2X2 U820 ( .A(n1092), .B(n1179), .Y(n1094) );
  OAI21X1 U821 ( .A0(n991), .A1(n147), .B0(n148), .Y(n1113) );
  XOR2X1TH U822 ( .A(n1140), .B(n1054), .Y(n778) );
  NOR2XLTH U823 ( .A(n1058), .B(n1188), .Y(n464) );
  NAND2X2TH U824 ( .A(n949), .B(n950), .Y(n740) );
  ADDFXLTH U825 ( .A(n332), .B(n468), .CI(n575), .CO(n327), .S(n328) );
  NOR2XLTH U826 ( .A(n1057), .B(n1191), .Y(n468) );
  INVX4TH U827 ( .A(n1141), .Y(n1175) );
  BUFX5 U828 ( .A(b[9]), .Y(n1133) );
  BUFX10 U829 ( .A(n784), .Y(n1146) );
  ADDFXL U830 ( .A(n282), .B(n293), .CI(n280), .CO(n277), .S(n278) );
  NAND3X2TH U831 ( .A(n883), .B(n884), .C(n885), .Y(n336) );
  BUFX8 U832 ( .A(b[11]), .Y(n1074) );
  NAND2X5TH U833 ( .A(n1108), .B(n95), .Y(n93) );
  CLKNAND2X4 U834 ( .A(n987), .B(n127), .Y(n125) );
  OR2X4 U835 ( .A(n128), .B(n126), .Y(n987) );
  NOR2X2 U836 ( .A(n266), .B(n277), .Y(n102) );
  INVX4 U837 ( .A(n1143), .Y(n1171) );
  NAND2X1TH U838 ( .A(n1172), .B(n1089), .Y(n1091) );
  CLKBUFX8 U839 ( .A(a[13]), .Y(n1144) );
  XNOR2X1 U840 ( .A(n117), .B(n63), .Y(product_18_) );
  BUFX4 U841 ( .A(b[14]), .Y(n1136) );
  INVX3TH U842 ( .A(n1144), .Y(n1167) );
  INVX5 U843 ( .A(n1124), .Y(n781) );
  NAND2X2 U844 ( .A(n954), .B(n955), .Y(product_28_) );
  CLKNAND2X2 U845 ( .A(n1149), .B(n1161), .Y(n955) );
  NAND2X4TH U846 ( .A(n932), .B(n933), .Y(n1066) );
  XNOR2X1TH U847 ( .A(n1136), .B(n1138), .Y(n741) );
  CLKNAND2X2TH U848 ( .A(n932), .B(n933), .Y(n1105) );
  OAI22XL U849 ( .A0(n694), .A1(n1096), .B0(n1070), .B1(n785), .Y(n544) );
  XNOR2X2 U851 ( .A(n1134), .B(n1141), .Y(n694) );
  BUFX10 U852 ( .A(n513), .Y(n1067) );
  BUFX6 U853 ( .A(n529), .Y(n1068) );
  XOR2X8 U854 ( .A(n311), .B(n481), .Y(n916) );
  OAI22X2 U855 ( .A0(n781), .A1(n632), .B0(n631), .B1(n1066), .Y(n481) );
  OAI22X1 U856 ( .A0(n1073), .A1(n666), .B0(n665), .B1(n1103), .Y(n514) );
  ADDFHX4 U857 ( .A(n560), .B(n1067), .CI(n349), .CO(n346), .S(n347) );
  OAI22X2 U858 ( .A0(n1073), .A1(n665), .B0(n664), .B1(n1103), .Y(n513) );
  BUFX20 U859 ( .A(n1075), .Y(n1069) );
  OAI22XL U860 ( .A0(n785), .A1(n699), .B0(n698), .B1(n1095), .Y(n548) );
  XNOR2X1 U861 ( .A(n1141), .B(n1130), .Y(n698) );
  BUFX6 U862 ( .A(n695), .Y(n1070) );
  XNOR2XL U863 ( .A(n1133), .B(n1141), .Y(n695) );
  INVX2 U864 ( .A(n1056), .Y(n1191) );
  NAND2XL U865 ( .A(n1139), .B(n1056), .Y(n964) );
  XNOR2X1 U866 ( .A(n1138), .B(n1056), .Y(n754) );
  OAI22XL U867 ( .A0(n723), .A1(n796), .B0(n724), .B1(n1147), .Y(n575) );
  XNOR2X2 U868 ( .A(n1133), .B(n1140), .Y(n712) );
  ADDFHX2 U869 ( .A(n591), .B(n345), .CI(n356), .CO(n340), .S(n341) );
  OAI22XL U870 ( .A0(n740), .A1(n1069), .B0(n1179), .B1(n1125), .Y(n591) );
  NOR2X2 U871 ( .A(n736), .B(n796), .Y(n967) );
  OAI22X2 U872 ( .A0(n1147), .A1(n736), .B0(n735), .B1(n796), .Y(n587) );
  XOR2XL U873 ( .A(n96), .B(n58), .Y(product_23_) );
  NAND2X1 U874 ( .A(n365), .B(n376), .Y(n132) );
  NAND3X2 U875 ( .A(n1027), .B(n1028), .C(n1029), .Y(n376) );
  CLKNAND2X4 U876 ( .A(n1182), .B(n1179), .Y(n888) );
  CLKINVX8 U877 ( .A(n1138), .Y(n1179) );
  ADDFHX2 U878 ( .A(n384), .B(n515), .CI(n593), .CO(n370), .S(n371) );
  OAI22X1 U879 ( .A0(n1073), .A1(n667), .B0(n666), .B1(n1103), .Y(n515) );
  OAI22X4 U880 ( .A0(n781), .A1(n635), .B0(n634), .B1(n1066), .Y(n484) );
  OAI22XL U881 ( .A0(n781), .A1(n633), .B0(n632), .B1(n1066), .Y(n482) );
  XNOR2XL U882 ( .A(n85), .B(n55), .Y(product_26_) );
  XOR2XL U883 ( .A(n112), .B(n62), .Y(product_19_) );
  XOR2XL U884 ( .A(n104), .B(n60), .Y(product_21_) );
  XNOR2XL U885 ( .A(n101), .B(n59), .Y(product_22_) );
  NOR2BX1 U886 ( .AN(n1148), .B(n1059), .Y(n469) );
  NOR2X4 U887 ( .A(n1059), .B(n1190), .Y(n467) );
  OAI22X4 U888 ( .A0(n1062), .A1(n719), .B0(n718), .B1(n795), .Y(n569) );
  OAI22X1 U889 ( .A0(n724), .A1(n796), .B0(n725), .B1(n1147), .Y(n576) );
  XNOR2X1 U890 ( .A(n1132), .B(n1140), .Y(n713) );
  ADDFHX1 U891 ( .A(n423), .B(n551), .CI(n598), .CO(n420), .S(n421) );
  ADDFHX1 U892 ( .A(n404), .B(n595), .CI(n503), .CO(n392), .S(n393) );
  NAND2XL U893 ( .A(n571), .B(n444), .Y(n961) );
  XOR2X8 U894 ( .A(n959), .B(n571), .Y(n441) );
  OAI22X4 U895 ( .A0(n1062), .A1(n721), .B0(n720), .B1(n795), .Y(n571) );
  XNOR2X1 U896 ( .A(n1140), .B(n1129), .Y(n716) );
  BUFX20 U897 ( .A(b[5]), .Y(n1129) );
  INVX20 U898 ( .A(b[12]), .Y(n1071) );
  CLKINVX40 U899 ( .A(n1071), .Y(n1072) );
  OAI22X2TH U900 ( .A0(n1147), .A1(n738), .B0(n737), .B1(n796), .Y(n589) );
  INVX2 U901 ( .A(n1137), .Y(n1180) );
  OAI22X2 U902 ( .A0(n729), .A1(n796), .B0(n730), .B1(n1147), .Y(n581) );
  ADDFHX1 U903 ( .A(n299), .B(n286), .CI(n297), .CO(n281), .S(n282) );
  CLKNAND2X2 U904 ( .A(n606), .B(n455), .Y(n182) );
  CLKNAND2X2TH U905 ( .A(n874), .B(n875), .Y(n720) );
  NAND2XLTH U906 ( .A(n1140), .B(n1128), .Y(n1085) );
  NOR2BXLTH U907 ( .AN(n1148), .B(n793), .Y(n536) );
  NOR2X2TH U908 ( .A(n904), .B(n868), .Y(n160) );
  ADDFX2TH U909 ( .A(n429), .B(n432), .CI(n427), .CO(n424), .S(n425) );
  XNOR2X1TH U910 ( .A(n1142), .B(n1128), .Y(n683) );
  ADDFXLTH U911 ( .A(n533), .B(n596), .CI(n405), .CO(n402), .S(n403) );
  INVX6 U912 ( .A(n1119), .Y(n796) );
  INVX2TH U913 ( .A(n1140), .Y(n1083) );
  INVXLTH U914 ( .A(n1128), .Y(n1084) );
  XOR2X3 U915 ( .A(n916), .B(n309), .Y(n294) );
  NAND3X2 U916 ( .A(n894), .B(n895), .C(n896), .Y(n253) );
  ADDFX1 U917 ( .A(n326), .B(n338), .CI(n324), .CO(n321), .S(n322) );
  NOR2X4TH U918 ( .A(n351), .B(n353), .Y(n126) );
  NAND2X2TH U919 ( .A(n351), .B(n353), .Y(n127) );
  BUFX12TH U920 ( .A(a[11]), .Y(n1143) );
  INVXLTH U921 ( .A(n1072), .Y(n1092) );
  XOR2X2TH U922 ( .A(n120), .B(n64), .Y(product_17_) );
  XOR2X1TH U923 ( .A(n72), .B(n52), .Y(product_29_) );
  BUFX8 U924 ( .A(a[1]), .Y(n1138) );
  NAND2X8 U925 ( .A(n775), .B(n1103), .Y(n1073) );
  NAND2X8 U926 ( .A(n774), .B(n791), .Y(n1077) );
  NAND2X6 U927 ( .A(n1081), .B(n1082), .Y(n746) );
  CLKNAND2X4 U928 ( .A(n1080), .B(n1179), .Y(n1082) );
  XNOR2XL U929 ( .A(n1128), .B(n1138), .Y(n751) );
  XNOR2X4 U930 ( .A(n1141), .B(n1128), .Y(n700) );
  BUFX20 U931 ( .A(b[4]), .Y(n1128) );
  OAI22XL U932 ( .A0(n727), .A1(n796), .B0(n728), .B1(n1147), .Y(n579) );
  NAND2BXL U933 ( .AN(n1148), .B(n1138), .Y(n756) );
  NAND2BXLTH U934 ( .AN(n1148), .B(n1139), .Y(n739) );
  NOR2BX4 U935 ( .AN(n1148), .B(n795), .Y(n572) );
  NOR2BXLTH U936 ( .AN(n1148), .B(n1095), .Y(n554) );
  BUFX12 U937 ( .A(n1060), .Y(n1148) );
  CLKNAND2X4 U938 ( .A(n1177), .B(n1191), .Y(n965) );
  CLKNAND2X4 U939 ( .A(n1186), .B(n1177), .Y(n1088) );
  CLKNAND2X2 U940 ( .A(n1177), .B(n1189), .Y(n881) );
  CLKNAND2X4 U941 ( .A(n1185), .B(n1177), .Y(n1039) );
  AND2X4 U942 ( .A(n1183), .B(n1177), .Y(n1104) );
  INVX3 U943 ( .A(n1139), .Y(n1177) );
  AO21XL U944 ( .A0(n1069), .A1(n1125), .B0(n1179), .Y(n319) );
  NAND2X1 U945 ( .A(n1180), .B(n1179), .Y(n950) );
  XOR2X3 U946 ( .A(n258), .B(n256), .Y(n893) );
  ADDFHX2 U947 ( .A(n260), .B(n478), .CI(n269), .CO(n255), .S(n256) );
  NAND2XL U948 ( .A(n1137), .B(n1138), .Y(n949) );
  XNOR2X4 U949 ( .A(n1137), .B(n1139), .Y(n723) );
  XNOR2X1 U950 ( .A(n1137), .B(n1141), .Y(n689) );
  XNOR2XL U951 ( .A(n1137), .B(n1142), .Y(n672) );
  XNOR2X1 U952 ( .A(n1128), .B(n1139), .Y(n734) );
  XNOR2X1 U953 ( .A(n1129), .B(n1139), .Y(n733) );
  NAND2X4 U954 ( .A(n1038), .B(n1039), .Y(n730) );
  XNOR2X1 U955 ( .A(n1133), .B(n1139), .Y(n729) );
  OAI22X1 U956 ( .A0(n746), .A1(n1125), .B0(n747), .B1(n1069), .Y(n598) );
  NAND2XL U957 ( .A(n1072), .B(n1138), .Y(n1093) );
  XNOR2XL U958 ( .A(n1072), .B(n1140), .Y(n709) );
  XNOR2XL U959 ( .A(n1072), .B(n1141), .Y(n692) );
  ADDFHX4 U960 ( .A(n581), .B(n407), .CI(n414), .CO(n404), .S(n405) );
  AND2X4 U961 ( .A(n565), .B(n549), .Y(n929) );
  OAI22X1 U962 ( .A0(n785), .A1(n700), .B0(n699), .B1(n1095), .Y(n549) );
  XNOR2X2 U963 ( .A(n125), .B(n65), .Y(product_16_) );
  CLKBUFX40 U964 ( .A(a[5]), .Y(n1140) );
  XOR2X1 U965 ( .A(n128), .B(n66), .Y(product_15_) );
  OAI22X2 U966 ( .A0(n741), .A1(n1125), .B0(n742), .B1(n1069), .Y(n593) );
  OAI22XL U967 ( .A0(n742), .A1(n1125), .B0(n743), .B1(n1069), .Y(n594) );
  CLKNAND2X2TH U968 ( .A(n887), .B(n888), .Y(n742) );
  NAND2XL U969 ( .A(n1131), .B(n1140), .Y(n1041) );
  NAND2X2 U970 ( .A(n1131), .B(n1139), .Y(n1087) );
  XNOR2X4 U971 ( .A(n1141), .B(n1131), .Y(n697) );
  XNOR2X4 U972 ( .A(n1131), .B(n1138), .Y(n748) );
  ADDHX4TH U973 ( .A(n604), .B(n589), .CO(n446), .S(n447) );
  ADDFHX1TH U974 ( .A(n586), .B(n442), .CI(n601), .CO(n438), .S(n439) );
  OAI22X2TH U975 ( .A0(n1055), .A1(n1125), .B0(n750), .B1(n1069), .Y(n601) );
  CLKNAND2X4 U976 ( .A(n117), .B(n866), .Y(n1106) );
  CLKAND2X2 U977 ( .A(n545), .B(n1068), .Y(n930) );
  XOR2X4TH U978 ( .A(n882), .B(n352), .Y(n337) );
  OR2X2 U979 ( .A(n278), .B(n291), .Y(n864) );
  OR2X4 U980 ( .A(n96), .B(n94), .Y(n1108) );
  NAND2X3 U981 ( .A(n939), .B(n940), .Y(n725) );
  NAND2X3 U982 ( .A(n779), .B(n796), .Y(n787) );
  CLKNAND2X2 U983 ( .A(n977), .B(n978), .Y(n777) );
  CLKNAND2X2 U984 ( .A(n1141), .B(n1176), .Y(n977) );
  NAND2X6 U985 ( .A(n983), .B(n103), .Y(n101) );
  INVX3 U986 ( .A(n110), .Y(n1150) );
  BUFX16 U987 ( .A(a[15]), .Y(n1145) );
  XNOR2X1TH U988 ( .A(n1127), .B(n1138), .Y(n752) );
  NOR2XLTH U989 ( .A(n1147), .B(n737), .Y(n966) );
  NOR2X1TH U990 ( .A(n605), .B(n590), .Y(n179) );
  XNOR2X1TH U991 ( .A(n1129), .B(n1138), .Y(n750) );
  NAND2X1 U992 ( .A(n1063), .B(n1159), .Y(n871) );
  CLKNAND2X2TH U993 ( .A(n1085), .B(n1086), .Y(n717) );
  NAND2X1TH U995 ( .A(n1083), .B(n1084), .Y(n1086) );
  NAND3X1TH U996 ( .A(n960), .B(n961), .C(n962), .Y(n440) );
  XNOR2X1TH U997 ( .A(n1141), .B(n1056), .Y(n703) );
  ADDFX1TH U998 ( .A(n566), .B(n422), .CI(n582), .CO(n414), .S(n415) );
  OAI22X1TH U999 ( .A0(n1146), .A1(n681), .B0(n680), .B1(n793), .Y(n529) );
  ADDFHXLTH U1000 ( .A(n519), .B(n420), .CI(n534), .CO(n410), .S(n411) );
  OAI22XLTH U1001 ( .A0(n1146), .A1(n686), .B0(n685), .B1(n793), .Y(n534) );
  OAI21X4TH U1002 ( .A0(n990), .A1(n155), .B0(n156), .Y(n1116) );
  NAND2XLTH U1003 ( .A(n425), .B(n430), .Y(n156) );
  NOR2XLTH U1004 ( .A(n425), .B(n430), .Y(n155) );
  OR2X1TH U1005 ( .A(n417), .B(n419), .Y(n1117) );
  OAI22XLTH U1006 ( .A0(n1146), .A1(n683), .B0(n682), .B1(n793), .Y(n531) );
  CLKNAND2X2TH U1007 ( .A(n876), .B(n877), .Y(n693) );
  NAND2XLTH U1008 ( .A(n1074), .B(n1141), .Y(n876) );
  INVXLTH U1009 ( .A(n319), .Y(n1156) );
  AND2XLTH U1010 ( .A(n1034), .B(n1035), .Y(n1019) );
  NAND2XLTH U1011 ( .A(n1136), .B(n1175), .Y(n1034) );
  NAND2XLTH U1012 ( .A(n1181), .B(n1141), .Y(n1035) );
  ADDFHXLTH U1013 ( .A(n303), .B(n1173), .CI(n509), .CO(n287), .S(n288) );
  INVXLTH U1014 ( .A(n289), .Y(n1173) );
  OAI22XLTH U1015 ( .A0(n1073), .A1(n661), .B0(n660), .B1(n1103), .Y(n509) );
  XNOR2X1TH U1016 ( .A(n1136), .B(n1140), .Y(n707) );
  ADDFXL U1017 ( .A(n512), .B(n334), .CI(n559), .CO(n331), .S(n332) );
  OAI22XLTH U1018 ( .A0(n708), .A1(n795), .B0(n709), .B1(n1062), .Y(n559) );
  NAND2XLTH U1019 ( .A(n902), .B(n903), .Y(n532) );
  OR2XLTH U1020 ( .A(n683), .B(n793), .Y(n903) );
  ADDFX1 U1021 ( .A(n510), .B(n304), .CI(n541), .CO(n301), .S(n302) );
  OAI22XLTH U1022 ( .A0(n691), .A1(n1096), .B0(n692), .B1(n785), .Y(n541) );
  NAND2X2TH U1023 ( .A(n969), .B(n970), .Y(n780) );
  ADDFX1TH U1024 ( .A(n517), .B(n395), .CI(n402), .CO(n390), .S(n391) );
  ADDFX1TH U1025 ( .A(n394), .B(n594), .CI(n392), .CO(n380), .S(n381) );
  AOI21X6TH U1026 ( .A0(n1113), .A1(n1114), .B0(n1115), .Y(n992) );
  OAI22XLTH U1027 ( .A0(n1077), .A1(n1167), .B0(n654), .B1(n791), .Y(n449) );
  NOR2BXLTH U1028 ( .AN(n1061), .B(n1105), .Y(n486) );
  ADDFX1 U1029 ( .A(n372), .B(n500), .CI(n370), .CO(n356), .S(n357) );
  OAI22XLTH U1030 ( .A0(n1077), .A1(n651), .B0(n650), .B1(n791), .Y(n500) );
  ADDFHX4TH U1031 ( .A(n592), .B(n359), .CI(n368), .CO(n354), .S(n355) );
  OAI22X1TH U1032 ( .A0(n740), .A1(n1125), .B0(n741), .B1(n1069), .Y(n592) );
  ADDFX1TH U1033 ( .A(n467), .B(n316), .CI(n574), .CO(n311), .S(n312) );
  ADDFHXLTH U1034 ( .A(n537), .B(n263), .CI(n507), .CO(n251), .S(n252) );
  OAI22XLTH U1035 ( .A0(n657), .A1(n1103), .B0(n1073), .B1(n658), .Y(n507) );
  NOR2X3TH U1036 ( .A(n292), .B(n305), .Y(n110) );
  CLKNAND2X2TH U1037 ( .A(n306), .B(n321), .Y(n116) );
  NAND2XLTH U1038 ( .A(n1153), .B(n127), .Y(n66) );
  XNOR2X1TH U1039 ( .A(n93), .B(n57), .Y(product_24_) );
  INVX2TH U1040 ( .A(n1074), .Y(n1183) );
  NAND2X1TH U1041 ( .A(a[10]), .B(n1142), .Y(n1090) );
  XOR2X1TH U1042 ( .A(n88), .B(n56), .Y(product_25_) );
  INVXLTH U1043 ( .A(n86), .Y(n1157) );
  INVXLTH U1044 ( .A(n77), .Y(n1149) );
  XOR2X1TH U1045 ( .A(n80), .B(n54), .Y(product_27_) );
  AND2X1TH U1046 ( .A(n773), .B(n1105), .Y(n1124) );
  XOR2XLTH U1047 ( .A(n1145), .B(n1079), .Y(n773) );
  XOR2X1TH U1048 ( .A(n1097), .B(n51), .Y(product_30_) );
  OA21X4TH U1049 ( .A0(n72), .A1(n70), .B0(n71), .Y(n1097) );
  XNOR2X1TH U1050 ( .A(n1135), .B(n1141), .Y(n691) );
  OAI22X1TH U1051 ( .A0(n1073), .A1(n660), .B0(n659), .B1(n1103), .Y(n508) );
  OAI22X1 U1052 ( .A0(n1073), .A1(n659), .B0(n658), .B1(n1103), .Y(n263) );
  NAND2X4 U1053 ( .A(n1167), .B(a[12]), .Y(n958) );
  CLKNAND2X4 U1054 ( .A(n1165), .B(n1167), .Y(n933) );
  OR2X6 U1055 ( .A(n898), .B(n899), .Y(n547) );
  NAND2XL U1056 ( .A(n339), .B(n341), .Y(n885) );
  ADDFHX4 U1057 ( .A(n343), .B(n484), .CI(n354), .CO(n338), .S(n339) );
  BUFX16 U1059 ( .A(a[9]), .Y(n1142) );
  INVX4 U1060 ( .A(n1142), .Y(n1089) );
  OR2X8 U1061 ( .A(n112), .B(n110), .Y(n1112) );
  NAND3X4 U1062 ( .A(n890), .B(n891), .C(n892), .Y(n299) );
  OAI22XL U1063 ( .A0(n1077), .A1(n649), .B0(n648), .B1(n791), .Y(n498) );
  CLKXOR2X2 U1064 ( .A(a[12]), .B(n1143), .Y(n1120) );
  OAI22X2 U1065 ( .A0(n725), .A1(n796), .B0(n726), .B1(n1147), .Y(n577) );
  OA21X4 U1066 ( .A0(n992), .A1(n139), .B0(n140), .Y(n136) );
  AND2X8 U1067 ( .A(n1107), .B(n92), .Y(n88) );
  XOR2X4 U1068 ( .A(n341), .B(n339), .Y(n882) );
  ADDFHX4 U1069 ( .A(n485), .B(n355), .CI(n364), .CO(n350), .S(n351) );
  OAI22X4 U1070 ( .A0(n712), .A1(n795), .B0(n713), .B1(n1062), .Y(n563) );
  AOI21X4 U1071 ( .A0(n1116), .A1(n1117), .B0(n1118), .Y(n991) );
  OAI22XL U1072 ( .A0(n1146), .A1(n682), .B0(n681), .B1(n793), .Y(n530) );
  CLKNAND2X2TH U1073 ( .A(n906), .B(n907), .Y(n682) );
  XNOR2X1 U1074 ( .A(n1134), .B(n1140), .Y(n711) );
  NAND2XL U1075 ( .A(n77), .B(n53), .Y(n954) );
  NAND2X5 U1076 ( .A(n1030), .B(n79), .Y(n77) );
  ADDFHX2 U1077 ( .A(n561), .B(n363), .CI(n374), .CO(n360), .S(n361) );
  XOR2X1 U1078 ( .A(n545), .B(n1068), .Y(n363) );
  ADDFX4 U1079 ( .A(n603), .B(n572), .CI(n588), .CO(n444), .S(n445) );
  OAI22XL U1080 ( .A0(n751), .A1(n1125), .B0(n752), .B1(n1069), .Y(n603) );
  OAI22XL U1081 ( .A0(n745), .A1(n1125), .B0(n746), .B1(n1069), .Y(n597) );
  ADDHX4 U1082 ( .A(n587), .B(n602), .CO(n442), .S(n443) );
  OAI22XL U1083 ( .A0(n750), .A1(n1125), .B0(n751), .B1(n1069), .Y(n602) );
  NAND2X8 U1084 ( .A(n936), .B(n937), .Y(n728) );
  CLKNAND2X4 U1085 ( .A(n1184), .B(n1177), .Y(n937) );
  NAND2XL U1086 ( .A(n1079), .B(n1144), .Y(n932) );
  BUFX6 U1087 ( .A(a[14]), .Y(n1079) );
  NOR2X6 U1088 ( .A(n322), .B(n336), .Y(n118) );
  OR2X4 U1089 ( .A(n337), .B(n350), .Y(n1049) );
  CLKNAND2X2 U1090 ( .A(n900), .B(n901), .Y(n452) );
  ADDFHX2TH U1091 ( .A(n451), .B(n421), .CI(n424), .CO(n416), .S(n417) );
  NAND2X3TH U1092 ( .A(n964), .B(n965), .Y(n737) );
  NOR2X2 U1093 ( .A(n441), .B(n453), .Y(n166) );
  CLKNAND2X2 U1094 ( .A(n1132), .B(n1139), .Y(n1038) );
  BUFX10 U1096 ( .A(b[3]), .Y(n1127) );
  INVX20 U1097 ( .A(n1102), .Y(n785) );
  AND2X6 U1098 ( .A(n777), .B(n1095), .Y(n1102) );
  NAND2X3 U1099 ( .A(n109), .B(n864), .Y(n1111) );
  CLKNAND2X2 U1100 ( .A(n926), .B(n84), .Y(n55) );
  XNOR2XLTH U1101 ( .A(n1138), .B(n1060), .Y(n755) );
  AND2XLTH U1102 ( .A(n605), .B(n590), .Y(n1020) );
  NAND2BXLTH U1103 ( .AN(n1148), .B(n1140), .Y(n722) );
  NAND2XLTH U1104 ( .A(n1140), .B(n1056), .Y(n874) );
  INVXLTH U1105 ( .A(n1063), .Y(n1178) );
  ADDFHXLTH U1106 ( .A(n600), .B(n435), .CI(n438), .CO(n432), .S(n433) );
  OAI22XLTH U1107 ( .A0(n748), .A1(n1125), .B0(n1055), .B1(n1069), .Y(n600) );
  CLKNAND2X2 U1108 ( .A(n871), .B(n872), .Y(n435) );
  ADDFHXLTH U1109 ( .A(n584), .B(n568), .CI(n928), .CO(n428), .S(n429) );
  AND2XLTH U1110 ( .A(n1063), .B(n569), .Y(n928) );
  OAI22X1TH U1111 ( .A0(n747), .A1(n1125), .B0(n748), .B1(n1069), .Y(n599) );
  XNOR2X1TH U1112 ( .A(n1142), .B(n1056), .Y(n686) );
  NOR2X2 U1113 ( .A(n437), .B(n440), .Y(n163) );
  NOR2XLTH U1114 ( .A(n431), .B(n433), .Y(n158) );
  NAND2XLTH U1115 ( .A(n431), .B(n433), .Y(n159) );
  ADDHXLTH U1116 ( .A(n547), .B(n563), .CO(n386), .S(n387) );
  OAI22X1TH U1117 ( .A0(n1070), .A1(n1095), .B0(n785), .B1(n696), .Y(n545) );
  ADDFX1TH U1118 ( .A(n550), .B(n597), .CI(n415), .CO(n412), .S(n413) );
  OAI22XLTH U1119 ( .A0(n785), .A1(n701), .B0(n700), .B1(n1095), .Y(n550) );
  OR2XLTH U1120 ( .A(n1146), .B(n684), .Y(n902) );
  ADDFHXLTH U1121 ( .A(n546), .B(n386), .CI(n562), .CO(n374), .S(n375) );
  OAI22XLTH U1122 ( .A0(n785), .A1(n697), .B0(n696), .B1(n1096), .Y(n546) );
  ADDFHXLTH U1123 ( .A(n319), .B(n573), .CI(n525), .CO(n303), .S(n304) );
  OAI22XLTH U1124 ( .A0(n676), .A1(n793), .B0(n1146), .B1(n677), .Y(n525) );
  NAND2XLTH U1125 ( .A(n1135), .B(n1139), .Y(n939) );
  NAND2XLTH U1126 ( .A(n1182), .B(n1177), .Y(n940) );
  OAI22XLTH U1127 ( .A0(n710), .A1(n795), .B0(n711), .B1(n1062), .Y(n561) );
  ADDFHXLTH U1129 ( .A(n544), .B(n528), .CI(n930), .CO(n348), .S(n349) );
  OAI22XLTH U1130 ( .A0(n1146), .A1(n680), .B0(n679), .B1(n793), .Y(n528) );
  NAND2XLTH U1131 ( .A(n1135), .B(n1138), .Y(n887) );
  NOR2BXLTH U1132 ( .AN(n1148), .B(n791), .Y(n503) );
  NAND2XLTH U1133 ( .A(n911), .B(n912), .Y(n533) );
  OR2XLTH U1134 ( .A(n1146), .B(n685), .Y(n911) );
  OR2XLTH U1135 ( .A(n399), .B(n401), .Y(n1114) );
  AND2XLTH U1136 ( .A(n399), .B(n401), .Y(n1115) );
  ADDFHXLTH U1137 ( .A(n530), .B(n578), .CI(n375), .CO(n372), .S(n373) );
  OAI22XLTH U1138 ( .A0(n726), .A1(n796), .B0(n727), .B1(n1147), .Y(n578) );
  XNOR2X1TH U1139 ( .A(n1144), .B(n1127), .Y(n650) );
  OAI22XLTH U1140 ( .A0(n692), .A1(n1096), .B0(n693), .B1(n785), .Y(n542) );
  OAI22XLTH U1141 ( .A0(n1146), .A1(n678), .B0(n677), .B1(n793), .Y(n526) );
  OAI22XLTH U1142 ( .A0(n706), .A1(n795), .B0(n707), .B1(n1062), .Y(n557) );
  CLKINVX4TH U1143 ( .A(a[0]), .Y(n1158) );
  ADDFHXLTH U1144 ( .A(n347), .B(n358), .CI(n469), .CO(n342), .S(n343) );
  OAI22XLTH U1145 ( .A0(n707), .A1(n795), .B0(n708), .B1(n1062), .Y(n558) );
  NAND2XLTH U1146 ( .A(n389), .B(n398), .Y(n140) );
  NOR2XLTH U1147 ( .A(n389), .B(n398), .Y(n139) );
  NAND2BXLTH U1148 ( .AN(n1061), .B(n1144), .Y(n654) );
  ADDFHXLTH U1149 ( .A(n373), .B(n486), .CI(n382), .CO(n368), .S(n369) );
  ADDFHXLTH U1150 ( .A(n482), .B(n312), .CI(n325), .CO(n307), .S(n308) );
  CLKINVX1TH U1151 ( .A(n1132), .Y(n1185) );
  CLKAND2X4TH U1152 ( .A(n938), .B(n135), .Y(n993) );
  CLKNAND2X2 U1153 ( .A(n377), .B(n379), .Y(n135) );
  OR2X4TH U1154 ( .A(n136), .B(n134), .Y(n938) );
  NOR2X3 U1155 ( .A(n377), .B(n379), .Y(n134) );
  XNOR2XLTH U1156 ( .A(n1145), .B(n1061), .Y(n636) );
  ADDFHXLTH U1157 ( .A(n310), .B(n323), .CI(n308), .CO(n305), .S(n306) );
  NAND2BXLTH U1158 ( .AN(n1101), .B(n793), .Y(n784) );
  AND2X6TH U1159 ( .A(n1106), .B(n116), .Y(n112) );
  INVXLTH U1160 ( .A(n1134), .Y(n1184) );
  NOR2X1TH U1161 ( .A(n233), .B(n226), .Y(n86) );
  NAND2XLTH U1162 ( .A(n1151), .B(n119), .Y(n64) );
  INVXLTH U1163 ( .A(n118), .Y(n1151) );
  NAND2XLTH U1164 ( .A(n1143), .B(n1172), .Y(n946) );
  OAI22X1TH U1165 ( .A0(n1077), .A1(n640), .B0(n639), .B1(n791), .Y(n223) );
  ADDFHXLTH U1166 ( .A(n231), .B(n222), .CI(n474), .CO(n219), .S(n220) );
  OAI22XLTH U1167 ( .A0(n781), .A1(n625), .B0(n624), .B1(n1066), .Y(n474) );
  OR2X1TH U1168 ( .A(n225), .B(n218), .Y(n926) );
  INVXLTH U1169 ( .A(n1079), .Y(n1165) );
  NAND2XLTH U1170 ( .A(n1162), .B(n79), .Y(n54) );
  NAND2XLTH U1171 ( .A(n994), .B(n68), .Y(n51) );
  NAND2XLTH U1172 ( .A(n199), .B(n201), .Y(n68) );
  NOR2X2TH U1173 ( .A(n244), .B(n253), .Y(n94) );
  XNOR2XL U1174 ( .A(n1139), .B(n1061), .Y(n738) );
  OAI22X1TH U1175 ( .A0(n730), .A1(n796), .B0(n731), .B1(n1147), .Y(n582) );
  AND2XLTH U1176 ( .A(n1074), .B(n1139), .Y(n1078) );
  INVXLTH U1177 ( .A(n1133), .Y(n1080) );
  XNOR2X1TH U1178 ( .A(n1145), .B(n1056), .Y(n635) );
  OAI22X1TH U1179 ( .A0(n1062), .A1(n1083), .B0(n722), .B1(n795), .Y(n453) );
  XNOR2X1TH U1180 ( .A(n1136), .B(n1139), .Y(n724) );
  NAND2XLTH U1181 ( .A(n481), .B(n311), .Y(n919) );
  AND2X8 U1182 ( .A(n1110), .B(n84), .Y(n80) );
  OR2X8 U1183 ( .A(n104), .B(n102), .Y(n983) );
  OAI22XL U1184 ( .A0(n1146), .A1(n687), .B0(n686), .B1(n793), .Y(n535) );
  OAI22XL U1185 ( .A0(n1146), .A1(n679), .B0(n678), .B1(n793), .Y(n527) );
  OAI22X4 U1186 ( .A0(n1062), .A1(n717), .B0(n716), .B1(n795), .Y(n567) );
  XNOR2X1 U1187 ( .A(n1132), .B(n1138), .Y(n747) );
  OA21X4 U1188 ( .A0(n988), .A1(n171), .B0(n172), .Y(n1099) );
  NOR2BX1 U1189 ( .AN(n1061), .B(n796), .Y(n590) );
  OAI22X4 U1190 ( .A0(n1069), .A1(n754), .B0(n753), .B1(n1125), .Y(n605) );
  OAI22X2 U1191 ( .A0(n752), .A1(n1125), .B0(n1069), .B1(n753), .Y(n604) );
  ADDFHX4 U1192 ( .A(n270), .B(n279), .CI(n268), .CO(n265), .S(n266) );
  NAND3X4 U1193 ( .A(n908), .B(n909), .C(n910), .Y(n279) );
  OAI22XLTH U1194 ( .A0(n713), .A1(n795), .B0(n714), .B1(n1062), .Y(n564) );
  OR2X6 U1195 ( .A(n1078), .B(n1104), .Y(n727) );
  NAND2BX1 U1196 ( .AN(n1148), .B(n1145), .Y(n637) );
  XNOR2X1 U1197 ( .A(n1074), .B(n1142), .Y(n676) );
  CLKNAND2X4 U1198 ( .A(n254), .B(n265), .Y(n100) );
  OR2X6 U1199 ( .A(n254), .B(n265), .Y(n865) );
  CLKXOR2X2TH U1200 ( .A(n893), .B(n267), .Y(n254) );
  XOR2X8 U1201 ( .A(n444), .B(n443), .Y(n959) );
  XNOR2X4 U1202 ( .A(n1134), .B(n1142), .Y(n677) );
  NAND2X3 U1203 ( .A(n93), .B(n925), .Y(n1107) );
  ADDFHX2TH U1204 ( .A(n396), .B(n516), .CI(n385), .CO(n382), .S(n383) );
  OAI22X2 U1205 ( .A0(n1073), .A1(n668), .B0(n667), .B1(n1103), .Y(n516) );
  OAI22X1TH U1206 ( .A0(n656), .A1(n1103), .B0(n657), .B1(n1073), .Y(n241) );
  CLKNAND2X2 U1207 ( .A(n225), .B(n218), .Y(n84) );
  OA21X2TH U1208 ( .A0(n160), .A1(n158), .B0(n159), .Y(n990) );
  ADDFHX1TH U1209 ( .A(n428), .B(n426), .CI(n535), .CO(n418), .S(n419) );
  CLKNAND2X2 U1210 ( .A(n256), .B(n258), .Y(n896) );
  CLKNAND2X2 U1211 ( .A(n267), .B(n256), .Y(n894) );
  OAI22X1TH U1212 ( .A0(n675), .A1(n793), .B0(n676), .B1(n1146), .Y(n289) );
  CLKNAND2X4 U1213 ( .A(n1087), .B(n1088), .Y(n731) );
  CLKNAND2X2 U1214 ( .A(n266), .B(n277), .Y(n103) );
  CLKNAND2X2 U1215 ( .A(n278), .B(n291), .Y(n108) );
  NOR2XLTH U1216 ( .A(n179), .B(n182), .Y(n1031) );
  OA21XLTH U1217 ( .A0(n174), .A1(n176), .B0(n175), .Y(n988) );
  NAND2XLTH U1218 ( .A(n447), .B(n1065), .Y(n175) );
  NOR2XLTH U1219 ( .A(n447), .B(n1065), .Y(n174) );
  NOR2XLTH U1220 ( .A(n1031), .B(n1020), .Y(n176) );
  NOR2XLTH U1221 ( .A(n445), .B(n446), .Y(n171) );
  OR2XLTH U1222 ( .A(n966), .B(n967), .Y(n588) );
  XNOR2XLTH U1223 ( .A(n1140), .B(n1061), .Y(n721) );
  NAND2XLTH U1224 ( .A(n1139), .B(n1127), .Y(n880) );
  NAND2XLTH U1225 ( .A(n445), .B(n446), .Y(n172) );
  NAND2XLTH U1226 ( .A(n443), .B(n444), .Y(n962) );
  ADDFHXLTH U1227 ( .A(n554), .B(n570), .CI(n439), .CO(n436), .S(n437) );
  OR2XLTH U1228 ( .A(n785), .B(n1175), .Y(n900) );
  ADDHX1TH U1229 ( .A(n567), .B(n583), .CO(n422), .S(n423) );
  NOR2X1TH U1230 ( .A(n989), .B(n163), .Y(n904) );
  NOR2X2TH U1231 ( .A(n897), .B(n867), .Y(n989) );
  AND2XLTH U1232 ( .A(n441), .B(n453), .Y(n867) );
  AND2XLTH U1233 ( .A(n437), .B(n440), .Y(n868) );
  XNOR2X1TH U1234 ( .A(n1141), .B(n1127), .Y(n701) );
  NOR2XLTH U1235 ( .A(n697), .B(n1095), .Y(n899) );
  ADDFHXLTH U1236 ( .A(n413), .B(n418), .CI(n411), .CO(n408), .S(n409) );
  INVXLTH U1237 ( .A(a[6]), .Y(n1176) );
  NAND2XLTH U1238 ( .A(n1175), .B(a[6]), .Y(n978) );
  ADDFHXLTH U1239 ( .A(n555), .B(n289), .CI(n508), .CO(n275), .S(n276) );
  AND2X1TH U1240 ( .A(n417), .B(n419), .Y(n1118) );
  NOR2XLTH U1241 ( .A(n409), .B(n416), .Y(n147) );
  NAND2XLTH U1242 ( .A(n409), .B(n416), .Y(n148) );
  ADDFHX2TH U1243 ( .A(n412), .B(n410), .CI(n518), .CO(n400), .S(n401) );
  XNOR2XLTH U1244 ( .A(n1144), .B(n1061), .Y(n653) );
  ADDFHXLTH U1245 ( .A(n315), .B(n466), .CI(n557), .CO(n297), .S(n298) );
  NAND2XLTH U1246 ( .A(n1021), .B(n1022), .Y(n510) );
  ADDFHXLTH U1247 ( .A(n540), .B(n495), .CI(n288), .CO(n285), .S(n286) );
  OAI22XLTH U1248 ( .A0(n1019), .A1(n1096), .B0(n691), .B1(n785), .Y(n540) );
  ADDFHXLTH U1249 ( .A(n524), .B(n276), .CI(n494), .CO(n273), .S(n274) );
  OAI22XLTH U1250 ( .A0(n674), .A1(n793), .B0(n675), .B1(n1146), .Y(n524) );
  OAI22XLTH U1251 ( .A0(n1077), .A1(n645), .B0(n644), .B1(n791), .Y(n494) );
  ADDFHXLTH U1252 ( .A(n287), .B(n464), .CI(n539), .CO(n271), .S(n272) );
  OAI22XLTH U1253 ( .A0(n689), .A1(n1096), .B0(n1019), .B1(n785), .Y(n539) );
  ADDFHXLTH U1254 ( .A(n493), .B(n463), .CI(n538), .CO(n259), .S(n260) );
  OAI22XLTH U1255 ( .A0(n689), .A1(n785), .B0(n1175), .B1(n1096), .Y(n538) );
  OAI22XLTH U1256 ( .A0(n1077), .A1(n644), .B0(n643), .B1(n791), .Y(n493) );
  ADDFHXLTH U1257 ( .A(n1169), .B(n523), .CI(n275), .CO(n261), .S(n262) );
  OAI22XLTH U1258 ( .A0(n673), .A1(n793), .B0(n674), .B1(n1146), .Y(n523) );
  INVXLTH U1259 ( .A(n263), .Y(n1169) );
  ADDFHXLTH U1260 ( .A(n344), .B(n330), .CI(n342), .CO(n325), .S(n326) );
  ADDFHXLTH U1261 ( .A(n328), .B(n483), .CI(n340), .CO(n323), .S(n324) );
  ADDFX1TH U1262 ( .A(n329), .B(n314), .CI(n327), .CO(n309), .S(n310) );
  OAI22XLTH U1263 ( .A0(n723), .A1(n1147), .B0(n1177), .B1(n796), .Y(n574) );
  NAND2XLTH U1264 ( .A(n302), .B(n317), .Y(n891) );
  ADDFX1TH U1265 ( .A(n301), .B(n465), .CI(n556), .CO(n283), .S(n284) );
  OAI22XLTH U1266 ( .A0(n706), .A1(n1062), .B0(n1083), .B1(n795), .Y(n556) );
  NOR2XLTH U1267 ( .A(n1058), .B(n1084), .Y(n465) );
  OAI22X1TH U1268 ( .A0(n781), .A1(n631), .B0(n630), .B1(n1066), .Y(n480) );
  ADDFHXLTH U1269 ( .A(n274), .B(n285), .CI(n283), .CO(n269), .S(n270) );
  ADDFX1TH U1270 ( .A(n272), .B(n479), .CI(n281), .CO(n267), .S(n268) );
  OAI22XLTH U1271 ( .A0(n781), .A1(n630), .B0(n629), .B1(n1066), .Y(n479) );
  ADDFX1TH U1273 ( .A(n262), .B(n273), .CI(n271), .CO(n257), .S(n258) );
  OAI22XLTH U1274 ( .A0(n781), .A1(n629), .B0(n628), .B1(n1066), .Y(n478) );
  XNOR2X1TH U1275 ( .A(n1135), .B(n1143), .Y(n657) );
  XNOR2X1TH U1276 ( .A(n1144), .B(n1074), .Y(n642) );
  ADDFHXLTH U1277 ( .A(n492), .B(n252), .CI(n462), .CO(n249), .S(n250) );
  NOR2XLTH U1278 ( .A(n1059), .B(n1186), .Y(n462) );
  ADDFHXLTH U1279 ( .A(n259), .B(n477), .CI(n257), .CO(n245), .S(n246) );
  OAI22XLTH U1280 ( .A0(n781), .A1(n628), .B0(n627), .B1(n1066), .Y(n477) );
  ADDFHXLTH U1282 ( .A(n522), .B(n261), .CI(n250), .CO(n247), .S(n248) );
  OAI22XLTH U1283 ( .A0(n672), .A1(n793), .B0(n673), .B1(n1146), .Y(n522) );
  NAND2XLTH U1284 ( .A(n381), .B(n390), .Y(n1029) );
  NAND2XLTH U1285 ( .A(n388), .B(n381), .Y(n1027) );
  NAND2XLTH U1286 ( .A(n388), .B(n390), .Y(n1028) );
  NAND2XLTH U1287 ( .A(n352), .B(n339), .Y(n883) );
  ADDFHXLTH U1288 ( .A(n296), .B(n307), .CI(n294), .CO(n291), .S(n292) );
  NAND2XLTH U1289 ( .A(n480), .B(n284), .Y(n910) );
  NAND2XLTH U1290 ( .A(n295), .B(n284), .Y(n909) );
  ADDFHXLTH U1291 ( .A(n248), .B(n255), .CI(n246), .CO(n243), .S(n244) );
  ADDFHXLTH U1292 ( .A(n1170), .B(n251), .CI(n491), .CO(n239), .S(n240) );
  OAI22XLTH U1293 ( .A0(n1077), .A1(n642), .B0(n641), .B1(n791), .Y(n491) );
  INVXLTH U1294 ( .A(n241), .Y(n1170) );
  ADDFHXLTH U1295 ( .A(n461), .B(n521), .CI(n240), .CO(n237), .S(n238) );
  OAI22XLTH U1296 ( .A0(n672), .A1(n1146), .B0(n1089), .B1(n793), .Y(n521) );
  NOR2XLTH U1297 ( .A(n1058), .B(n1185), .Y(n461) );
  ADDFHXLTH U1298 ( .A(n249), .B(n476), .CI(n238), .CO(n235), .S(n236) );
  OAI22XLTH U1299 ( .A0(n781), .A1(n627), .B0(n626), .B1(n1066), .Y(n476) );
  ADDFHXLTH U1300 ( .A(n247), .B(n236), .CI(n245), .CO(n233), .S(n234) );
  OR2X1TH U1301 ( .A(n306), .B(n321), .Y(n866) );
  NAND2XLTH U1302 ( .A(n234), .B(n243), .Y(n92) );
  OR2XLTH U1303 ( .A(n234), .B(n243), .Y(n925) );
  NAND2X1TH U1304 ( .A(n244), .B(n253), .Y(n95) );
  XNOR2X1TH U1305 ( .A(n1144), .B(n1135), .Y(n640) );
  NAND2XLTH U1306 ( .A(n1171), .B(a[10]), .Y(n947) );
  ADDFHXLTH U1307 ( .A(n520), .B(n241), .CI(n490), .CO(n231), .S(n232) );
  OAI22XLTH U1308 ( .A0(n1077), .A1(n641), .B0(n640), .B1(n791), .Y(n490) );
  ADDFHXLTH U1309 ( .A(n460), .B(n506), .CI(n232), .CO(n229), .S(n230) );
  NOR2XLTH U1310 ( .A(n1059), .B(n1080), .Y(n460) );
  OAI22XLTH U1311 ( .A0(n655), .A1(n1103), .B0(n656), .B1(n1073), .Y(n506) );
  ADDFHXLTH U1312 ( .A(n239), .B(n475), .CI(n230), .CO(n227), .S(n228) );
  OAI22XLTH U1313 ( .A0(n781), .A1(n626), .B0(n625), .B1(n1066), .Y(n475) );
  ADDFHXLTH U1314 ( .A(n237), .B(n228), .CI(n235), .CO(n225), .S(n226) );
  NAND2XLTH U1315 ( .A(n866), .B(n116), .Y(n63) );
  INVXLTH U1316 ( .A(n102), .Y(n1155) );
  NAND2XLTH U1317 ( .A(n1150), .B(n111), .Y(n62) );
  NAND2XLTH U1318 ( .A(n925), .B(n92), .Y(n57) );
  NAND2XLTH U1319 ( .A(n864), .B(n108), .Y(n61) );
  NAND2XLTH U1320 ( .A(n865), .B(n100), .Y(n59) );
  NAND2XLTH U1321 ( .A(n1154), .B(n95), .Y(n58) );
  INVXLTH U1322 ( .A(n94), .Y(n1154) );
  NAND2XLTH U1323 ( .A(n1157), .B(n87), .Y(n56) );
  ADDFHXLTH U1324 ( .A(n229), .B(n227), .CI(n220), .CO(n217), .S(n218) );
  ADDFHXLTH U1325 ( .A(n1166), .B(n459), .CI(n505), .CO(n221), .S(n222) );
  NOR2XLTH U1326 ( .A(n1058), .B(n1184), .Y(n459) );
  INVXLTH U1327 ( .A(n223), .Y(n1166) );
  NAND2XLTH U1328 ( .A(n927), .B(n76), .Y(n53) );
  ADDFHXLTH U1329 ( .A(n504), .B(n223), .CI(n458), .CO(n215), .S(n216) );
  NOR2XLTH U1330 ( .A(n1059), .B(n1183), .Y(n458) );
  ADDFHXLTH U1331 ( .A(n473), .B(n214), .CI(n219), .CO(n211), .S(n212) );
  OAI22XLTH U1332 ( .A0(n781), .A1(n624), .B0(n623), .B1(n1066), .Y(n473) );
  NOR2XLTH U1333 ( .A(n217), .B(n212), .Y(n78) );
  NAND2XLTH U1334 ( .A(n217), .B(n212), .Y(n79) );
  ADDFHXLTH U1335 ( .A(n489), .B(n216), .CI(n221), .CO(n213), .S(n214) );
  OAI22XLTH U1337 ( .A0(n638), .A1(n791), .B0(n1077), .B1(n639), .Y(n489) );
  ADDFHXLTH U1338 ( .A(n488), .B(n1163), .CI(n215), .CO(n207), .S(n208) );
  OAI22XLTH U1339 ( .A0(n638), .A1(n1077), .B0(n1167), .B1(n791), .Y(n488) );
  INVXLTH U1340 ( .A(n209), .Y(n1163) );
  XNOR2X1TH U1341 ( .A(n1145), .B(n1137), .Y(n621) );
  ADDFHXLTH U1342 ( .A(n487), .B(n209), .CI(n457), .CO(n203), .S(n204) );
  NOR2XLTH U1343 ( .A(n1059), .B(n1182), .Y(n457) );
  OR2XLTH U1344 ( .A(n211), .B(n206), .Y(n927) );
  NAND2XLTH U1345 ( .A(n211), .B(n206), .Y(n76) );
  ADDFHXLTH U1346 ( .A(n472), .B(n208), .CI(n213), .CO(n205), .S(n206) );
  OAI22XLTH U1347 ( .A0(n781), .A1(n623), .B0(n622), .B1(n1066), .Y(n472) );
  NAND2XLTH U1348 ( .A(n1160), .B(n71), .Y(n52) );
  INVXLTH U1349 ( .A(n70), .Y(n1160) );
  ADDFHXLTH U1350 ( .A(n204), .B(n471), .CI(n207), .CO(n201), .S(n202) );
  OAI22XLTH U1351 ( .A0(n781), .A1(n622), .B0(n621), .B1(n1066), .Y(n471) );
  XOR3XLTH U1352 ( .A(n456), .B(n203), .C(n1100), .Y(n199) );
  NOR2XLTH U1353 ( .A(n1058), .B(n1181), .Y(n456) );
  OR2XLTH U1354 ( .A(n199), .B(n201), .Y(n994) );
  NAND2XLTH U1355 ( .A(n1133), .B(n1138), .Y(n1081) );
  OAI22XLTH U1356 ( .A0(n1062), .A1(n718), .B0(n717), .B1(n795), .Y(n568) );
  OAI22X2 U1357 ( .A0(n731), .A1(n796), .B0(n732), .B1(n1147), .Y(n583) );
  OAI22XLTH U1358 ( .A0(n1073), .A1(n1171), .B0(n671), .B1(n1103), .Y(n450) );
  OAI22XL U1359 ( .A0(n1073), .A1(n663), .B0(n662), .B1(n1103), .Y(n511) );
  OAI22XLTH U1360 ( .A0(n655), .A1(n1073), .B0(n1171), .B1(n1103), .Y(n505) );
  XOR2X3 U1361 ( .A(n1064), .B(n1138), .Y(n1119) );
  XNOR2X1TH U1362 ( .A(n1141), .B(n1129), .Y(n699) );
  CLKINVX40 U1363 ( .A(n1122), .Y(n793) );
  AND2X8 U1364 ( .A(n1174), .B(n1175), .Y(n1123) );
  CLKXOR2X4 U1365 ( .A(n1054), .B(n1139), .Y(n1121) );
  CLKINVX24 U1366 ( .A(n1121), .Y(n795) );
  OR2X4 U1367 ( .A(n80), .B(n78), .Y(n1030) );
  NAND2XLTH U1368 ( .A(n233), .B(n226), .Y(n87) );
  NAND2X8 U1369 ( .A(n101), .B(n865), .Y(n1109) );
  NAND2XLTH U1370 ( .A(n205), .B(n202), .Y(n71) );
  OR2XLTH U1371 ( .A(n684), .B(n793), .Y(n912) );
  NOR2BX8 U1372 ( .AN(n1024), .B(n1123), .Y(n1122) );
  CLKINVX1TH U1373 ( .A(n1127), .Y(n1189) );
  BUFX20 U1374 ( .A(n787), .Y(n1147) );
  XNOR2X1TH U1375 ( .A(n1140), .B(n1127), .Y(n718) );
  INVXLTH U1376 ( .A(a[12]), .Y(n1168) );
  XNOR2X1TH U1377 ( .A(n1135), .B(n1140), .Y(n708) );
  INVXLTH U1378 ( .A(n78), .Y(n1162) );
  NAND2XLTH U1379 ( .A(n267), .B(n258), .Y(n895) );
  NOR2XLTH U1380 ( .A(n205), .B(n202), .Y(n70) );
  ADDFHX2 U1381 ( .A(n357), .B(n366), .CI(n448), .CO(n352), .S(n353) );
  OAI22XLTH U1382 ( .A0(n1077), .A1(n646), .B0(n645), .B1(n791), .Y(n495) );
  OAI22XLTH U1383 ( .A0(n1077), .A1(n643), .B0(n642), .B1(n791), .Y(n492) );
  OA22XLTH U1384 ( .A0(n781), .A1(n621), .B0(n1059), .B1(n1066), .Y(n1100) );
  XNOR2X1 U1385 ( .A(n1134), .B(n1138), .Y(n745) );
  INVX12 U1386 ( .A(n1120), .Y(n791) );
  XOR2XL U1387 ( .A(n1139), .B(n1064), .Y(n779) );
  XNOR2X4 U1388 ( .A(a[6]), .B(n1140), .Y(n1095) );
  XNOR2X4 U1389 ( .A(a[6]), .B(n1140), .Y(n1096) );
  AOI21BX4 U1390 ( .A0(n77), .A1(n927), .B0N(n76), .Y(n72) );
  AND2X6 U1391 ( .A(n1109), .B(n100), .Y(n96) );
  AND2X6 U1392 ( .A(n1111), .B(n108), .Y(n104) );
  NAND2XLTH U1393 ( .A(n1155), .B(n103), .Y(n60) );
  INVXLTH U1394 ( .A(n1049), .Y(n1152) );
  INVXLTH U1395 ( .A(n569), .Y(n1159) );
  NAND2XLTH U1396 ( .A(n352), .B(n341), .Y(n884) );
  NAND2XLTH U1397 ( .A(n1178), .B(n569), .Y(n872) );
  NAND2XLTH U1398 ( .A(n295), .B(n480), .Y(n908) );
  NAND2XLTH U1399 ( .A(n309), .B(n481), .Y(n917) );
  NAND2XLTH U1400 ( .A(n309), .B(n311), .Y(n918) );
  OAI22XLTH U1401 ( .A0(n1062), .A1(n720), .B0(n719), .B1(n795), .Y(n570) );
  NOR2XLTH U1402 ( .A(n1058), .B(n1187), .Y(n463) );
  XNOR2XLTH U1403 ( .A(n1143), .B(n1061), .Y(n670) );
  INVXLTH U1404 ( .A(a[10]), .Y(n1172) );
  NAND2XLTH U1406 ( .A(n1142), .B(n1127), .Y(n914) );
  XNOR2X1TH U1407 ( .A(n1132), .B(n1141), .Y(n696) );
  XNOR2X1TH U1408 ( .A(n1074), .B(n1140), .Y(n710) );
  XNOR2X1TH U1409 ( .A(n1142), .B(n1132), .Y(n679) );
  XNOR2X1TH U1410 ( .A(n1142), .B(n1131), .Y(n680) );
  XNOR2X1TH U1411 ( .A(n1142), .B(n1130), .Y(n681) );
  XNOR2X1TH U1412 ( .A(n1143), .B(n1130), .Y(n664) );
  XNOR2X1TH U1413 ( .A(n1143), .B(n1129), .Y(n665) );
  XNOR2X1TH U1414 ( .A(n1144), .B(n1126), .Y(n651) );
  XNOR2X1TH U1415 ( .A(n1143), .B(n1056), .Y(n669) );
  XNOR2X1TH U1416 ( .A(n1143), .B(n1128), .Y(n666) );
  XNOR2X1TH U1417 ( .A(n1144), .B(n1128), .Y(n649) );
  XNOR2X1TH U1418 ( .A(n1145), .B(n1126), .Y(n634) );
  XNOR2X1TH U1419 ( .A(n1144), .B(n1056), .Y(n652) );
  XNOR2X1TH U1420 ( .A(n1143), .B(n1127), .Y(n667) );
  INVXLTH U1421 ( .A(n1126), .Y(n1190) );
  NAND2XLTH U1422 ( .A(n1142), .B(n1129), .Y(n906) );
  NAND2XLTH U1423 ( .A(n1134), .B(n1139), .Y(n936) );
  XNOR2X1TH U1424 ( .A(n1143), .B(n1131), .Y(n663) );
  XNOR2X1TH U1425 ( .A(n1144), .B(n1131), .Y(n646) );
  XNOR2X1TH U1426 ( .A(n1145), .B(n1129), .Y(n631) );
  XNOR2X1TH U1427 ( .A(n1142), .B(n1133), .Y(n678) );
  XNOR2X1TH U1428 ( .A(n1144), .B(n1130), .Y(n647) );
  XNOR2X1TH U1429 ( .A(n1145), .B(n1130), .Y(n630) );
  XNOR2X1TH U1430 ( .A(n1145), .B(n1128), .Y(n632) );
  XNOR2X1TH U1431 ( .A(n1144), .B(n1129), .Y(n648) );
  XNOR2X1TH U1432 ( .A(n1143), .B(n1132), .Y(n662) );
  XNOR2X1TH U1433 ( .A(n1143), .B(n1133), .Y(n661) );
  XNOR2X1TH U1434 ( .A(n1145), .B(n1127), .Y(n633) );
  XNOR2XLTH U1435 ( .A(n1141), .B(n1061), .Y(n704) );
  INVXLTH U1436 ( .A(n1136), .Y(n1181) );
  INVXLTH U1437 ( .A(n1129), .Y(n1188) );
  NAND2BXLTH U1438 ( .AN(n1061), .B(n1141), .Y(n705) );
  XNOR2X1TH U1439 ( .A(n1136), .B(n1142), .Y(n673) );
  XNOR2X1TH U1440 ( .A(n1136), .B(n1143), .Y(n656) );
  XNOR2X1TH U1441 ( .A(n1072), .B(n1143), .Y(n658) );
  XNOR2X1TH U1442 ( .A(n1143), .B(n1134), .Y(n660) );
  XNOR2X1TH U1443 ( .A(n1144), .B(n1134), .Y(n643) );
  XNOR2X1TH U1444 ( .A(n1145), .B(n1132), .Y(n628) );
  XNOR2X1TH U1445 ( .A(n1144), .B(n1132), .Y(n645) );
  XNOR2X1TH U1446 ( .A(n1145), .B(n1131), .Y(n629) );
  XNOR2X1TH U1447 ( .A(n1145), .B(n1133), .Y(n627) );
  XNOR2X1TH U1448 ( .A(n1144), .B(n1133), .Y(n644) );
  XNOR2X1TH U1449 ( .A(n1135), .B(n1142), .Y(n674) );
  XNOR2X1TH U1450 ( .A(n1137), .B(n1143), .Y(n655) );
  XNOR2X1TH U1451 ( .A(n1136), .B(n1144), .Y(n639) );
  XNOR2X1TH U1452 ( .A(n1145), .B(n1074), .Y(n625) );
  XNOR2X1TH U1453 ( .A(n1145), .B(n1134), .Y(n626) );
  XNOR2X1TH U1454 ( .A(n1144), .B(n1072), .Y(n641) );
  NOR2XLTH U1455 ( .A(n1058), .B(n1092), .Y(n209) );
  XNOR2X1TH U1456 ( .A(n1137), .B(n1144), .Y(n638) );
  XNOR2X1TH U1457 ( .A(n1145), .B(n1136), .Y(n622) );
  XNOR2X1TH U1458 ( .A(n1145), .B(n1072), .Y(n624) );
  XNOR2X1TH U1459 ( .A(n1145), .B(n1135), .Y(n623) );
  INVXLTH U1460 ( .A(n1130), .Y(n1187) );
  AO21XLTH U1461 ( .A0(n1062), .A1(n795), .B0(n1083), .Y(n555) );
  ADDFX1 U1462 ( .A(n333), .B(n511), .CI(n318), .CO(n315), .S(n316) );
  XOR3XL U1463 ( .A(n295), .B(n480), .C(n284), .Y(n280) );
  ADDFX1 U1464 ( .A(n553), .B(n452), .CI(n436), .CO(n430), .S(n431) );
  OR2XLTH U1465 ( .A(n705), .B(n1095), .Y(n901) );
  ADDFX1 U1466 ( .A(n1156), .B(n527), .CI(n543), .CO(n333), .S(n334) );
  OR2XLTH U1467 ( .A(n661), .B(n1103), .Y(n1022) );
  OAI22XLTH U1468 ( .A0(n709), .A1(n795), .B0(n710), .B1(n1062), .Y(n560) );
  ADDFX1TH U1469 ( .A(n1156), .B(n526), .CI(n542), .CO(n317), .S(n318) );
  OR2XLTH U1470 ( .A(n1073), .B(n662), .Y(n1021) );
  AO21XLTH U1471 ( .A0(n785), .A1(n1096), .B0(n1175), .Y(n537) );
  AO21XLTH U1472 ( .A0(n1147), .A1(n796), .B0(n1177), .Y(n573) );
  AO21XLTH U1473 ( .A0(n1073), .A1(n1103), .B0(n1171), .Y(n504) );
  AO21XLTH U1474 ( .A0(n1146), .A1(n793), .B0(n1089), .Y(n520) );
  AO21XLTH U1475 ( .A0(n1077), .A1(n791), .B0(n1167), .Y(n487) );
  OAI22XLTH U1476 ( .A0(n1077), .A1(n653), .B0(n652), .B1(n791), .Y(n502) );
  NAND2XLTH U1477 ( .A(n1089), .B(n1189), .Y(n915) );
  NAND2XLTH U1479 ( .A(n1089), .B(n1188), .Y(n907) );
  NAND2XLTH U1480 ( .A(n1083), .B(n1191), .Y(n875) );
  ADDFX1 U1481 ( .A(n450), .B(n403), .CI(n408), .CO(n398), .S(n399) );
  NAND2XLTH U1482 ( .A(n1186), .B(n1083), .Y(n1042) );
  NAND2XLTH U1483 ( .A(n1183), .B(n1175), .Y(n877) );
  INVXL U1484 ( .A(n53), .Y(n1161) );
endmodule


module multiplier_1 ( data1, data2, out );
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] out;
  wire   N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, abs_data2_15_, N87, N88, N89, N90, N91, N92, N93,
         N94, N95, N96, N97, N98, N99, N100, N101, N102, n7, n9, n10, n19, n20,
         n210, n220, n230, n240, n250, n260, n270, n280, n290, n320, n38, n1,
         n2, n3, n4, n5, n6, n11, n14, n17, n18, n300, n310, n330, n350, n360,
         n39, n40, n41, n44, n46, n50, n51, n52, n53, n540, n550, n560, n570,
         n600, n610, n640, n660, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165;
  wire   [15:0] abs_data1;
  wire   [30:15] abs_c;

  INVXL U51 ( .A(abs_c[27]), .Y(n4) );
  NOR2BX1 U98 ( .AN(N36), .B(n310), .Y(abs_data1[15]) );
  multiplier_1_DW01_inc_0 add_41 ( .A({n1, n2, n3, n4, n5, n6, n132, n11, n133, 
        n136, n14, n135, n137, n17, n18, n300}), .SUM({N102, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87}) );
  multiplier_1_DW01_inc_1 add_29 ( .A({n165, n50, n51, n52, n53, n540, n550, 
        n560, n570, n158, n157, n600, n610, n155, n154, n640}), .SUM({N69, N68, 
        N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54})
         );
  multiplier_1_DW01_inc_2 add_21 ( .A({n310, n330, n153, n350, n360, n150, n39, 
        n40, n41, n148, n147, n44, n146, n46, n145, n144}), .SUM({N36, N35, 
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21})
         );
  multiplier_1_DW_mult_uns_3 mult_36 ( .a({abs_data1[15:10], n660, 
        abs_data1[8:2], n19, abs_data1[0]}), .b({abs_data2_15_, n320, n10, 
        n270, n9, n7, n250, n240, n280, n260, n230, n290, n210, n220, n38, 
        n143}), .product_30_(abs_c[30]), .product_29_(abs_c[29]), 
        .product_28_(abs_c[28]), .product_27_(abs_c[27]), .product_26_(
        abs_c[26]), .product_25_(abs_c[25]), .product_24_(abs_c[24]), 
        .product_23_(abs_c[23]), .product_22_(abs_c[22]), .product_21_(
        abs_c[21]), .product_20_(abs_c[20]), .product_19_(abs_c[19]), 
        .product_18_(abs_c[18]), .product_17_(abs_c[17]), .product_16_(
        abs_c[16]), .product_15_(abs_c[15]) );
  AO2B2X2 U2 ( .B0(N92), .B1(n140), .A0(n134), .A1N(n139), .Y(out[5]) );
  OAI2B2XL U3 ( .A1N(N25), .A0(n310), .B0(n123), .B1(n44), .Y(abs_data1[4]) );
  INVX20 U4 ( .A(n123), .Y(n310) );
  OAI2B2X4 U5 ( .A1N(N63), .A0(n165), .B0(data2[15]), .B1(n161), .Y(n250) );
  BUFX6 U6 ( .A(abs_c[22]), .Y(n128) );
  BUFX6 U7 ( .A(n20), .Y(n143) );
  CLKBUFX40 U8 ( .A(data1[15]), .Y(n123) );
  INVX2TH U9 ( .A(data1[2]), .Y(n46) );
  INVX4TH U10 ( .A(data1[1]), .Y(n145) );
  CLKBUFX2TH U11 ( .A(abs_c[23]), .Y(n124) );
  CLKBUFX2TH U12 ( .A(abs_c[21]), .Y(n127) );
  CLKINVX1TH U13 ( .A(data1[7]), .Y(n41) );
  AO2B2X4 U14 ( .B0(N89), .B1(n140), .A0(abs_c[17]), .A1N(n139), .Y(out[2]) );
  INVX2 U15 ( .A(abs_c[17]), .Y(n17) );
  OAI2B2XL U16 ( .A1N(N35), .A0(n310), .B0(n123), .B1(n330), .Y(abs_data1[14])
         );
  BUFX6 U17 ( .A(abs_c[26]), .Y(n125) );
  BUFX6 U18 ( .A(abs_c[19]), .Y(n126) );
  INVX4 U19 ( .A(abs_c[24]), .Y(n132) );
  AO2B2X4 U20 ( .B0(N96), .B1(n141), .A0(abs_c[24]), .A1N(n139), .Y(out[9]) );
  AO2B2X4 U21 ( .B0(N101), .B1(n140), .A0(abs_c[29]), .A1N(n139), .Y(out[14])
         );
  INVX2 U22 ( .A(abs_c[29]), .Y(n2) );
  INVX2TH U23 ( .A(n127), .Y(n136) );
  CLKINVX1TH U24 ( .A(data1[6]), .Y(n148) );
  CLKINVX1TH U25 ( .A(data2[5]), .Y(n157) );
  CLKINVX1TH U26 ( .A(data1[5]), .Y(n147) );
  CLKINVX1TH U27 ( .A(data2[6]), .Y(n158) );
  AO2B2XLTH U28 ( .B0(N98), .B1(n141), .A0(n125), .A1N(n140), .Y(out[11]) );
  CLKINVX1TH U29 ( .A(data1[13]), .Y(n153) );
  CLKINVX1TH U30 ( .A(data1[9]), .Y(n39) );
  OAI2B2X4 U31 ( .A1N(data1[1]), .A0(n123), .B0(n138), .B1(n310), .Y(n19) );
  OAI2B2XL U32 ( .A1N(N23), .A0(n310), .B0(n123), .B1(n46), .Y(abs_data1[2])
         );
  OAI2B2X4 U33 ( .A1N(N31), .A0(n310), .B0(n123), .B1(n150), .Y(abs_data1[10])
         );
  CLKINVX40 U34 ( .A(data2[15]), .Y(n165) );
  OAI2B2X4 U35 ( .A1N(N58), .A0(n165), .B0(data2[15]), .B1(n156), .Y(n290) );
  OAI2B2XLTH U36 ( .A1N(N54), .A0(n165), .B0(data2[15]), .B1(n640), .Y(n20) );
  OAI2B2X4 U37 ( .A1N(N62), .A0(n165), .B0(data2[15]), .B1(n160), .Y(n240) );
  OAI2B2XLTH U38 ( .A1N(N56), .A0(n165), .B0(data2[15]), .B1(n155), .Y(n220)
         );
  INVX1TH U39 ( .A(data2[2]), .Y(n155) );
  INVX2TH U40 ( .A(data2[1]), .Y(n154) );
  BUFX6 U41 ( .A(abs_c[15]), .Y(n129) );
  OAI2B2X4 U42 ( .A1N(N67), .A0(n165), .B0(data2[15]), .B1(n164), .Y(n10) );
  CLKINVX3TH U43 ( .A(data2[0]), .Y(n640) );
  OAI2B2X4TH U44 ( .A1N(N29), .A0(n310), .B0(n123), .B1(n149), .Y(abs_data1[8]) );
  OAI2B2X4TH U45 ( .A1N(N30), .A0(n310), .B0(n123), .B1(n39), .Y(n660) );
  BUFX4 U46 ( .A(abs_c[20]), .Y(n134) );
  INVX2TH U47 ( .A(abs_c[16]), .Y(n18) );
  INVX2TH U48 ( .A(n129), .Y(n300) );
  INVXLTH U49 ( .A(n128), .Y(n133) );
  INVXLTH U50 ( .A(data2[13]), .Y(n164) );
  CLKBUFX2 U52 ( .A(abs_c[25]), .Y(n131) );
  NOR2BXLTH U53 ( .AN(N69), .B(n165), .Y(abs_data2_15_) );
  INVXLTH U54 ( .A(abs_c[28]), .Y(n3) );
  INVX1TH U55 ( .A(data1[3]), .Y(n146) );
  INVX1TH U56 ( .A(n126), .Y(n135) );
  XNOR2XLTH U57 ( .A(n310), .B(data2[15]), .Y(n130) );
  OAI2B2X4 U58 ( .A1N(N33), .A0(n310), .B0(n123), .B1(n152), .Y(abs_data1[12])
         );
  AO2B2X4 U59 ( .B0(N21), .B1(n123), .A0(n310), .A1N(n144), .Y(abs_data1[0])
         );
  OAI2B2X4 U60 ( .A1N(N26), .A0(n310), .B0(n123), .B1(n147), .Y(abs_data1[5])
         );
  OAI2B2X4 U61 ( .A1N(N28), .A0(n310), .B0(n123), .B1(n41), .Y(abs_data1[7])
         );
  OAI2B2X4 U62 ( .A1N(N55), .A0(n165), .B0(data2[15]), .B1(n154), .Y(n38) );
  AO2B2X1 U63 ( .B0(N88), .B1(n140), .A0(abs_c[16]), .A1N(n139), .Y(out[1]) );
  INVX6 U64 ( .A(abs_c[18]), .Y(n137) );
  OAI2B2X4TH U65 ( .A1N(N59), .A0(n165), .B0(data2[15]), .B1(n157), .Y(n230)
         );
  OAI2B2X4TH U66 ( .A1N(N57), .A0(n165), .B0(data2[15]), .B1(n610), .Y(n210)
         );
  INVXLTH U67 ( .A(data2[4]), .Y(n156) );
  INVXLTH U68 ( .A(data2[7]), .Y(n159) );
  INVXLTH U69 ( .A(data2[9]), .Y(n161) );
  OAI2B2X2TH U70 ( .A1N(N64), .A0(n165), .B0(data2[15]), .B1(n540), .Y(n7) );
  INVXLTH U71 ( .A(data2[11]), .Y(n162) );
  OAI2B2X4TH U72 ( .A1N(N66), .A0(n165), .B0(data2[15]), .B1(n163), .Y(n270)
         );
  INVXLTH U73 ( .A(data2[12]), .Y(n163) );
  INVXLTH U74 ( .A(n134), .Y(n14) );
  INVXLTH U75 ( .A(data1[14]), .Y(n330) );
  OAI2B2X4TH U76 ( .A1N(N32), .A0(n310), .B0(n123), .B1(n151), .Y(
        abs_data1[11]) );
  INVXLTH U77 ( .A(data1[11]), .Y(n151) );
  AO2B2XLTH U78 ( .B0(N91), .B1(n140), .A0(n126), .A1N(n139), .Y(out[4]) );
  AO2B2XLTH U79 ( .B0(N95), .B1(n141), .A0(n124), .A1N(n139), .Y(out[8]) );
  OAI2B2X4TH U80 ( .A1N(N68), .A0(n165), .B0(data2[15]), .B1(n50), .Y(n320) );
  INVXLTH U81 ( .A(n131), .Y(n6) );
  CLKINVX1TH U82 ( .A(data1[4]), .Y(n44) );
  AO2B2XLTH U83 ( .B0(N97), .B1(n141), .A0(n131), .A1N(n140), .Y(out[10]) );
  AO2B2XLTH U84 ( .B0(N93), .B1(n141), .A0(n127), .A1N(n139), .Y(out[6]) );
  AO2B2XLTH U85 ( .B0(N94), .B1(n141), .A0(n128), .A1N(n139), .Y(out[7]) );
  AO2B2XLTH U86 ( .B0(N90), .B1(n140), .A0(abs_c[18]), .A1N(n139), .Y(out[3])
         );
  OAI2B2X4 U87 ( .A1N(N61), .A0(n165), .B0(data2[15]), .B1(n159), .Y(n280) );
  OAI2B2X4 U88 ( .A1N(N65), .A0(n165), .B0(data2[15]), .B1(n162), .Y(n9) );
  INVX2TH U89 ( .A(n124), .Y(n11) );
  OAI2B2X4 U90 ( .A1N(N24), .A0(n310), .B0(n123), .B1(n146), .Y(abs_data1[3])
         );
  INVX1TH U91 ( .A(abs_c[30]), .Y(n1) );
  CLKINVX12TH U92 ( .A(data1[0]), .Y(n144) );
  INVXLTH U93 ( .A(data2[3]), .Y(n610) );
  INVXLTH U94 ( .A(data2[4]), .Y(n600) );
  INVXLTH U95 ( .A(data2[7]), .Y(n570) );
  INVXLTH U96 ( .A(data2[8]), .Y(n560) );
  INVXLTH U97 ( .A(data2[8]), .Y(n160) );
  INVXLTH U99 ( .A(data1[8]), .Y(n40) );
  INVXLTH U100 ( .A(data1[8]), .Y(n149) );
  INVXLTH U101 ( .A(data2[9]), .Y(n550) );
  INVXLTH U102 ( .A(data2[10]), .Y(n540) );
  INVXLTH U103 ( .A(data2[11]), .Y(n53) );
  INVXLTH U104 ( .A(data1[10]), .Y(n150) );
  INVXLTH U105 ( .A(data1[12]), .Y(n350) );
  INVXLTH U106 ( .A(data1[11]), .Y(n360) );
  INVXLTH U107 ( .A(data2[12]), .Y(n52) );
  INVXLTH U108 ( .A(data2[13]), .Y(n51) );
  CLKBUFX2TH U109 ( .A(n142), .Y(n141) );
  INVXLTH U110 ( .A(data2[14]), .Y(n50) );
  INVXLTH U111 ( .A(data1[12]), .Y(n152) );
  AO2B2XLTH U112 ( .B0(N87), .B1(n141), .A0(n129), .A1N(n140), .Y(out[0]) );
  AO2B2XLTH U113 ( .B0(N99), .B1(n140), .A0(abs_c[27]), .A1N(n140), .Y(out[12]) );
  AO2B2XLTH U114 ( .B0(N100), .B1(n140), .A0(abs_c[28]), .A1N(n139), .Y(
        out[13]) );
  INVXLTH U115 ( .A(n125), .Y(n5) );
  CLKBUFX1TH U116 ( .A(n130), .Y(n142) );
  BUFX3TH U117 ( .A(n142), .Y(n140) );
  CLKBUFX3TH U118 ( .A(n142), .Y(n139) );
  OAI2B2X4 U119 ( .A1N(N34), .A0(n310), .B0(n123), .B1(n153), .Y(abs_data1[13]) );
  INVX4 U120 ( .A(N22), .Y(n138) );
  OAI2BB2X4 U121 ( .B0(n1), .B1(n139), .A0N(N102), .A1N(n140), .Y(out[15]) );
  OAI2B2X4 U122 ( .A1N(N27), .A0(n310), .B0(n123), .B1(n148), .Y(abs_data1[6])
         );
  OAI2B2X1 U123 ( .A1N(N60), .A0(n165), .B0(data2[15]), .B1(n158), .Y(n260) );
endmodule


module multiplier_0_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;
  wire   n1, n2, n3;
  wire   [15:2] carry;

  ADDHX2 U1_1_5 ( .A(A[5]), .B(n1), .CO(carry[6]), .S(SUM[5]) );
  ADDHX4TH U1_1_3 ( .A(A[3]), .B(n2), .CO(carry[4]), .S(SUM[3]) );
  ADDHX2TH U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXLTH U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHX2TH U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXLTH U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXLTH U1_1_11 ( .A(A[11]), .B(n3), .CO(carry[12]), .S(SUM[11]) );
  ADDHX2 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX2TH U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXLTH U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  AND2X8 U1 ( .A(A[4]), .B(carry[4]), .Y(n1) );
  XOR2X2 U2 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  CLKAND2X4TH U3 ( .A(A[2]), .B(carry[2]), .Y(n2) );
  XOR2X1 U4 ( .A(A[10]), .B(carry[10]), .Y(SUM[10]) );
  XOR2XLTH U5 ( .A(A[4]), .B(carry[4]), .Y(SUM[4]) );
  AND2XLTH U6 ( .A(A[10]), .B(carry[10]), .Y(n3) );
  XOR2XLTH U7 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
  INVXLTH U8 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module multiplier_0_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  ADDHXLTH U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXLTH U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXLTH U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXLTH U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXLTH U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXLTH U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXLTH U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXLTH U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXLTH U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXLTH U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXLTH U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXLTH U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXLTH U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXLTH U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR2XLTH U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  INVXLTH U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module multiplier_0_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;
  wire   n3, n4, n5, n6, n8, n11, n12, n13, n14, n15, n16;
  wire   [14:2] carry;

  INVXL U13 ( .A(A[0]), .Y(SUM[0]) );
  ADDHX2TH U1_1_13 ( .A(A[13]), .B(n5), .CO(carry[14]), .S(SUM[13]) );
  ADDHXLTH U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXLTH U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXLTH U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXLTH U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXLTH U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXLTH U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHX4 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHX4 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_11 ( .A(A[11]), .B(n8), .CO(carry[12]), .S(SUM[11]) );
  ADDHX1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVXLTH U1 ( .A(A[10]), .Y(n16) );
  XOR2X3 U2 ( .A(A[12]), .B(carry[12]), .Y(SUM[12]) );
  XOR2X3 U3 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  AND2X6 U4 ( .A(A[10]), .B(carry[10]), .Y(n8) );
  NAND2X2TH U5 ( .A(n14), .B(A[15]), .Y(n4) );
  CLKNAND2X2TH U6 ( .A(n3), .B(n4), .Y(SUM[15]) );
  CLKNAND2X2 U7 ( .A(n11), .B(n12), .Y(SUM[10]) );
  AND2XLTH U8 ( .A(A[14]), .B(carry[14]), .Y(n6) );
  INVXLTH U9 ( .A(carry[10]), .Y(n13) );
  NAND2XLTH U10 ( .A(n16), .B(carry[10]), .Y(n12) );
  AND2X4 U11 ( .A(A[12]), .B(carry[12]), .Y(n5) );
  INVXLTH U12 ( .A(n6), .Y(n14) );
  NAND2XLTH U14 ( .A(n6), .B(n15), .Y(n3) );
  INVXLTH U15 ( .A(A[15]), .Y(n15) );
  NAND2XLTH U16 ( .A(A[10]), .B(n13), .Y(n11) );
endmodule


module multiplier_0_DW_mult_uns_3 ( a, b, product_30_, product_29_, 
        product_28_, product_27_, product_26_, product_25_, product_24_, 
        product_23_, product_22_, product_21_, product_20_, product_19_, 
        product_18_, product_17_, product_16_, product_15_ );
  input [15:0] a;
  input [15:0] b;
  output product_30_, product_29_, product_28_, product_27_, product_26_,
         product_25_, product_24_, product_23_, product_22_, product_21_,
         product_20_, product_19_, product_18_, product_17_, product_16_,
         product_15_;
  wire   n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n68, n69, n70, n71, n72, n76, n77, n79, n80, n84, n85, n87,
         n88, n92, n93, n95, n96, n100, n101, n102, n103, n104, n108, n109,
         n110, n111, n112, n116, n117, n118, n119, n120, n124, n125, n126,
         n127, n128, n131, n132, n134, n139, n140, n142, n144, n147, n148,
         n150, n152, n155, n156, n163, n164, n166, n167, n168, n171, n174,
         n175, n176, n179, n180, n182, n199, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n443, n444, n445, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n773, n774, n775, n776,
         n777, n778, n779, n780, n788, n790, n791, n792, n793, n794, n795,
         n796, n862, n863, n867, n868, n873, n874, n875, n876, n879, n880,
         n881, n882, n884, n885, n886, n887, n888, n889, n891, n892, n893,
         n894, n897, n898, n899, n900, n902, n903, n906, n907, n909, n910,
         n911, n912, n913, n914, n916, n917, n918, n919, n920, n923, n924,
         n925, n926, n927, n928, n929, n930, n932, n933, n935, n936, n937,
         n938, n939, n940, n941, n944, n947, n949, n950, n951, n952, n953,
         n954, n957, n958, n960, n961, n963, n964, n968, n969, n970, n972,
         n973, n975, n976, n985, n988, n994, n996, n997, n998, n999, n1001,
         n1012, n1013, n1014, n1017, n1018, n1020, n1021, n1022, n1023, n1025,
         n1026, n1028, n1029, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1044, n1045, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165;

  NOR2X2TH U891 ( .A(n365), .B(n376), .Y(n131) );
  NOR2X2 U715 ( .A(n399), .B(n408), .Y(n142) );
  NAND2X2 U902 ( .A(n881), .B(n882), .Y(n571) );
  NOR2BX1 U1261 ( .AN(n1124), .B(n794), .Y(n554) );
  OAI22X1 U1273 ( .A0(n661), .A1(n1052), .B0(n660), .B1(n792), .Y(n508) );
  NAND2X2 U890 ( .A(n1153), .B(n1165), .Y(n1026) );
  OAI22X1 U956 ( .A0(n735), .A1(n796), .B0(n736), .B1(n1050), .Y(n587) );
  NOR2X1 U1013 ( .A(n445), .B(n929), .Y(n171) );
  OAI22X1 U1041 ( .A0(n633), .A1(n790), .B0(n634), .B1(n1048), .Y(n479) );
  OAI22X1 U1062 ( .A0(n665), .A1(n792), .B0(n666), .B1(n1052), .Y(n513) );
  NAND2BX2 U1065 ( .AN(n1123), .B(n1107), .Y(n637) );
  NAND2X2 U1470 ( .A(n1150), .B(n1160), .Y(n973) );
  ADDFX1 U707 ( .A(n387), .B(n396), .CI(n394), .CO(n380), .S(n381) );
  XNOR2X1 U708 ( .A(n1118), .B(n1101), .Y(n727) );
  BUFX10 U709 ( .A(a[11]), .Y(n1118) );
  NOR2X6 U710 ( .A(n144), .B(n142), .Y(n941) );
  CLKNAND2X12 U711 ( .A(n944), .B(n95), .Y(n93) );
  NAND2X5 U712 ( .A(n1129), .B(n867), .Y(n944) );
  CLKNAND2X12 U713 ( .A(n1082), .B(n103), .Y(n101) );
  OR2X8 U714 ( .A(n104), .B(n102), .Y(n1082) );
  CLKNAND2X12 U716 ( .A(n1083), .B(n111), .Y(n109) );
  OR2X8 U717 ( .A(n112), .B(n110), .Y(n1083) );
  NOR2X4 U718 ( .A(n930), .B(n928), .Y(n997) );
  AND2X1 U719 ( .A(n417), .B(n424), .Y(n928) );
  NOR2X8 U720 ( .A(n152), .B(n150), .Y(n930) );
  BUFX12 U721 ( .A(a[2]), .Y(n1109) );
  NAND2X2 U722 ( .A(n1127), .B(n1058), .Y(n985) );
  OA21X2 U723 ( .A0(n179), .A1(n182), .B0(n180), .Y(n176) );
  NOR2XL U724 ( .A(n605), .B(n590), .Y(n179) );
  NAND2X2 U725 ( .A(n85), .B(n924), .Y(n1086) );
  CLKNAND2X8 U726 ( .A(n947), .B(n87), .Y(n85) );
  NAND2X4 U727 ( .A(n1065), .B(n1066), .Y(n605) );
  OAI22X1 U728 ( .A0(n740), .A1(n1099), .B0(n741), .B1(n788), .Y(n592) );
  NAND2X8 U729 ( .A(n957), .B(n958), .Y(n740) );
  OR2X2 U730 ( .A(n742), .B(n1099), .Y(n1034) );
  OAI22X1 U731 ( .A0(n742), .A1(n788), .B0(n741), .B1(n1099), .Y(n593) );
  CLKNAND2X4 U732 ( .A(n963), .B(n964), .Y(n742) );
  NOR2XL U733 ( .A(n409), .B(n416), .Y(n147) );
  ADDFHX4 U734 ( .A(n413), .B(n418), .CI(n411), .CO(n408), .S(n409) );
  XOR2XL U735 ( .A(n104), .B(n60), .Y(product_21_) );
  AND2X8 U736 ( .A(n988), .B(n108), .Y(n104) );
  ADDFHX4 U737 ( .A(n360), .B(n345), .CI(n591), .CO(n340), .S(n341) );
  OAI22XLTH U738 ( .A0(n740), .A1(n788), .B0(n1165), .B1(n1099), .Y(n591) );
  ADDFHX2 U739 ( .A(n480), .B(n576), .CI(n362), .CO(n344), .S(n345) );
  XOR2X1 U740 ( .A(n128), .B(n66), .Y(product_15_) );
  CLKNAND2X4 U741 ( .A(n863), .B(n116), .Y(n63) );
  CLKNAND2X2 U742 ( .A(n306), .B(n321), .Y(n116) );
  OAI22X2 U743 ( .A0(n729), .A1(n796), .B0(n730), .B1(n1050), .Y(n581) );
  OR2X2 U744 ( .A(n729), .B(n1050), .Y(n1040) );
  XNOR2X1 U745 ( .A(n1116), .B(n1101), .Y(n729) );
  NAND2X6 U746 ( .A(n1028), .B(n1029), .Y(n718) );
  NAND2X2 U747 ( .A(n606), .B(n455), .Y(n182) );
  OAI22X1TH U748 ( .A0(n755), .A1(n788), .B0(n754), .B1(n1099), .Y(n606) );
  CLKNAND2X4 U749 ( .A(n891), .B(n892), .Y(n682) );
  NOR2XL U750 ( .A(n1154), .B(n1156), .Y(n464) );
  CLKNAND2X4 U751 ( .A(n1154), .B(n1159), .Y(n894) );
  CLKNAND2X4 U752 ( .A(n1154), .B(n1163), .Y(n910) );
  INVX1 U753 ( .A(n1108), .Y(n1154) );
  BUFX20 U754 ( .A(a[12]), .Y(n1119) );
  CLKNAND2X4 U755 ( .A(n1125), .B(n62), .Y(n880) );
  INVX6 U756 ( .A(n62), .Y(n1133) );
  CLKNAND2X4 U757 ( .A(n1134), .B(n111), .Y(n62) );
  XNOR2X1 U758 ( .A(n1115), .B(n1102), .Y(n713) );
  BUFX12 U759 ( .A(a[8]), .Y(n1115) );
  BUFX10 U760 ( .A(n449), .Y(n1047) );
  CLKNAND2X4 U761 ( .A(n968), .B(n969), .Y(n741) );
  ADDFHX4 U762 ( .A(n326), .B(n338), .CI(n324), .CO(n321), .S(n322) );
  NAND3X2 U763 ( .A(n1037), .B(n1038), .C(n1039), .Y(n338) );
  CLKNAND2X2TH U764 ( .A(n322), .B(n336), .Y(n119) );
  NOR2X8 U765 ( .A(n322), .B(n336), .Y(n118) );
  NAND3X2 U766 ( .A(n952), .B(n953), .C(n954), .Y(n336) );
  ADDFHX2 U767 ( .A(n310), .B(n323), .CI(n308), .CO(n305), .S(n306) );
  NAND2X4 U768 ( .A(n437), .B(n440), .Y(n164) );
  NOR2X6 U769 ( .A(n437), .B(n440), .Y(n163) );
  CLKXOR2X2 U770 ( .A(n911), .B(n439), .Y(n437) );
  OR2X8 U771 ( .A(n120), .B(n118), .Y(n1084) );
  INVX6 U772 ( .A(n118), .Y(n1132) );
  XOR2XL U773 ( .A(n120), .B(n64), .Y(product_17_) );
  OR2X4 U774 ( .A(n337), .B(n350), .Y(n862) );
  NAND2X3 U775 ( .A(n337), .B(n350), .Y(n124) );
  NAND3X4 U776 ( .A(n938), .B(n939), .C(n940), .Y(n350) );
  OR2X8 U777 ( .A(n728), .B(n796), .Y(n1041) );
  OAI22X4 U778 ( .A0(n727), .A1(n796), .B0(n728), .B1(n1050), .Y(n579) );
  XNOR2X4 U779 ( .A(n1117), .B(n1101), .Y(n728) );
  XOR2X8 U780 ( .A(n951), .B(n339), .Y(n337) );
  XOR2X8 U781 ( .A(n1036), .B(n343), .Y(n339) );
  NAND2X4 U782 ( .A(n893), .B(n894), .Y(n686) );
  INVX2 U783 ( .A(n1112), .Y(n1149) );
  BUFX10 U784 ( .A(a[1]), .Y(n1108) );
  XOR2X1TH U785 ( .A(n80), .B(n54), .Y(product_27_) );
  AND2X1TH U786 ( .A(n453), .B(n602), .Y(n873) );
  CLKNAND2X4 U787 ( .A(n916), .B(n917), .Y(n701) );
  NAND2X2 U788 ( .A(n1152), .B(n1163), .Y(n917) );
  ADDFXLTH U789 ( .A(n309), .B(n307), .CI(n294), .CO(n291), .S(n292) );
  OAI22XLTH U790 ( .A0(n731), .A1(n1050), .B0(n730), .B1(n796), .Y(n582) );
  CLKBUFX6 U791 ( .A(a[5]), .Y(n1112) );
  BUFX10 U792 ( .A(a[4]), .Y(n1111) );
  BUFX3 U793 ( .A(a[0]), .Y(n1056) );
  BUFX5 U794 ( .A(a[9]), .Y(n1116) );
  INVX2 U795 ( .A(n1047), .Y(n1155) );
  CLKBUFX4 U796 ( .A(a[14]), .Y(n1121) );
  BUFX8TH U797 ( .A(n1056), .Y(n1123) );
  XOR2X4 U798 ( .A(n72), .B(n52), .Y(product_29_) );
  XNOR2X1TH U799 ( .A(n1122), .B(n1101), .Y(n723) );
  OAI22X1 U800 ( .A0(n725), .A1(n1050), .B0(n724), .B1(n796), .Y(n576) );
  OAI22X1TH U801 ( .A0(n725), .A1(n796), .B0(n726), .B1(n1050), .Y(n577) );
  ADDFX1TH U802 ( .A(n359), .B(n361), .CI(n370), .CO(n354), .S(n355) );
  NAND2X4TH U803 ( .A(n773), .B(n790), .Y(n1048) );
  NAND2X4TH U804 ( .A(n774), .B(n791), .Y(n1049) );
  XNOR2X1TH U805 ( .A(n1110), .B(n1100), .Y(n752) );
  NAND2X4 U806 ( .A(n779), .B(n796), .Y(n1050) );
  XNOR2XL U807 ( .A(n101), .B(n59), .Y(product_22_) );
  XNOR2XL U808 ( .A(n109), .B(n61), .Y(product_20_) );
  NAND2X5 U809 ( .A(n1074), .B(n71), .Y(n69) );
  OR2X6 U810 ( .A(n72), .B(n70), .Y(n1074) );
  CLKNAND2X4 U811 ( .A(n897), .B(n898), .Y(n731) );
  OR2X4 U812 ( .A(n750), .B(n1099), .Y(n1063) );
  CLKNAND2X8 U813 ( .A(n109), .B(n868), .Y(n988) );
  INVX2 U814 ( .A(n88), .Y(n1128) );
  CLKNAND2X4 U815 ( .A(n1025), .B(n1026), .Y(n753) );
  NAND2XLTH U816 ( .A(n1109), .B(n1100), .Y(n1025) );
  XNOR2X1TH U817 ( .A(n1108), .B(n1100), .Y(n754) );
  XNOR2X1TH U818 ( .A(n1108), .B(n1101), .Y(n737) );
  XNOR2X1TH U819 ( .A(n1111), .B(n1100), .Y(n751) );
  XOR2X1 U820 ( .A(n873), .B(n601), .Y(n911) );
  NAND2XLTH U821 ( .A(n972), .B(n973), .Y(n734) );
  ADDFXLTH U822 ( .A(n1151), .B(n508), .CI(n540), .CO(n287), .S(n288) );
  NAND2XLTH U823 ( .A(n439), .B(n601), .Y(n912) );
  ADDFXLTH U824 ( .A(n569), .B(n600), .CI(n553), .CO(n432), .S(n433) );
  ADDFXLTH U825 ( .A(n435), .B(n438), .CI(n433), .CO(n430), .S(n431) );
  ADDFXLTH U826 ( .A(n552), .B(n584), .CI(n434), .CO(n426), .S(n427) );
  NAND2X2TH U827 ( .A(n960), .B(n961), .Y(n744) );
  XNOR2X1 U828 ( .A(n1119), .B(n1100), .Y(n743) );
  XOR2XLTH U829 ( .A(n451), .B(n567), .Y(n423) );
  ADDFX1TH U830 ( .A(n421), .B(n426), .CI(n419), .CO(n416), .S(n417) );
  OR2XLTH U831 ( .A(n743), .B(n788), .Y(n1035) );
  ADDFXLTH U832 ( .A(n1013), .B(n415), .CI(n420), .CO(n410), .S(n411) );
  ADDFXLTH U833 ( .A(n414), .B(n412), .CI(n405), .CO(n400), .S(n401) );
  OAI22X1 U834 ( .A0(n654), .A1(n791), .B0(n1049), .B1(n1157), .Y(n449) );
  NAND2X1TH U835 ( .A(n975), .B(n976), .Y(n726) );
  AND2X6 U836 ( .A(n101), .B(n876), .Y(n1076) );
  ADDFXLTH U837 ( .A(n403), .B(n410), .CI(n401), .CO(n398), .S(n399) );
  ADDFXLTH U838 ( .A(n393), .B(n400), .CI(n391), .CO(n388), .S(n389) );
  ADDFXLTH U839 ( .A(n404), .B(n395), .CI(n402), .CO(n390), .S(n391) );
  OR2XLTH U840 ( .A(n1057), .B(n1081), .Y(n724) );
  OAI22XLTH U841 ( .A0(n637), .A1(n790), .B0(n1048), .B1(n1156), .Y(n448) );
  ADDFXLTH U842 ( .A(n381), .B(n390), .CI(n379), .CO(n376), .S(n377) );
  OAI22XLTH U843 ( .A0(n723), .A1(n1050), .B0(n796), .B1(n1160), .Y(n574) );
  NAND2X6 U844 ( .A(n1084), .B(n119), .Y(n117) );
  NAND2X2 U845 ( .A(n1142), .B(n1165), .Y(n969) );
  INVX2 U846 ( .A(n1121), .Y(n1142) );
  NAND2X2 U847 ( .A(n1070), .B(n1071), .Y(n755) );
  XNOR2X1 U848 ( .A(n1117), .B(n1103), .Y(n694) );
  BUFX20 U849 ( .A(a[10]), .Y(n1117) );
  NAND2XL U850 ( .A(n1122), .B(n1100), .Y(n957) );
  BUFX12 U851 ( .A(a[15]), .Y(n1122) );
  CLKNAND2X4 U852 ( .A(n1144), .B(n1164), .Y(n936) );
  INVXL U853 ( .A(n1119), .Y(n1144) );
  OAI22X1 U854 ( .A0(n731), .A1(n796), .B0(n732), .B1(n1050), .Y(n583) );
  AOI21X8 U855 ( .A0(n1087), .A1(n1088), .B0(n1089), .Y(n999) );
  OAI21X8 U856 ( .A0(n1001), .A1(n163), .B0(n164), .Y(n1087) );
  NAND2X4 U857 ( .A(n1047), .B(n1140), .Y(n1017) );
  OAI22XL U858 ( .A0(n723), .A1(n796), .B0(n724), .B1(n1050), .Y(n575) );
  OA21X4 U859 ( .A0(n997), .A1(n147), .B0(n148), .Y(n144) );
  XNOR2X1 U860 ( .A(n1120), .B(n1101), .Y(n725) );
  NOR2X1TH U861 ( .A(n377), .B(n388), .Y(n134) );
  CLKNAND2X4 U862 ( .A(n935), .B(n936), .Y(n709) );
  CLKNAND2X4 U863 ( .A(n1072), .B(n1073), .Y(n453) );
  XNOR2X1 U864 ( .A(n1108), .B(n1102), .Y(n720) );
  NAND2XL U865 ( .A(n1108), .B(n1104), .Y(n893) );
  XNOR2X1 U866 ( .A(n1108), .B(n1106), .Y(n652) );
  CLKNAND2X2 U867 ( .A(n601), .B(n873), .Y(n914) );
  NOR2X1 U868 ( .A(n417), .B(n424), .Y(n150) );
  XNOR2XL U869 ( .A(n117), .B(n63), .Y(product_18_) );
  NAND2X2TH U870 ( .A(n1141), .B(n1165), .Y(n958) );
  NAND2X5 U871 ( .A(n909), .B(n910), .Y(n703) );
  XOR2X8 U872 ( .A(n356), .B(n354), .Y(n1036) );
  OAI22X1 U873 ( .A0(n750), .A1(n788), .B0(n749), .B1(n1099), .Y(n601) );
  CLKNAND2X4 U874 ( .A(n906), .B(n907), .Y(n750) );
  NOR2X2 U875 ( .A(n1080), .B(n171), .Y(n918) );
  CLKNAND2X2 U876 ( .A(n447), .B(n589), .Y(n175) );
  CLKNAND2X2 U877 ( .A(n1111), .B(n1101), .Y(n972) );
  AND2X2 U878 ( .A(n431), .B(n436), .Y(n1089) );
  ADDFHX2TH U879 ( .A(n429), .B(n432), .CI(n427), .CO(n424), .S(n425) );
  NAND2X3 U880 ( .A(n949), .B(n950), .Y(n745) );
  INVX4TH U881 ( .A(n69), .Y(n1126) );
  NAND2X3 U882 ( .A(n1128), .B(n1014), .Y(n947) );
  XOR2X1TH U883 ( .A(n88), .B(n56), .Y(product_25_) );
  OAI21X8TH U884 ( .A0(n128), .A1(n126), .B0(n127), .Y(n125) );
  OAI22XLTH U885 ( .A0(n756), .A1(n1099), .B0(n788), .B1(n1165), .Y(n455) );
  OR2XLTH U886 ( .A(n754), .B(n788), .Y(n1065) );
  NOR2BXLTH U887 ( .AN(n1124), .B(n796), .Y(n590) );
  NAND2XLTH U888 ( .A(n1061), .B(n1062), .Y(n604) );
  NAND2XLTH U889 ( .A(n1059), .B(n1060), .Y(n454) );
  CLKXOR2X2 U892 ( .A(n454), .B(n604), .Y(n447) );
  NOR2X2TH U893 ( .A(n447), .B(n589), .Y(n174) );
  AND2X1TH U894 ( .A(n454), .B(n604), .Y(n929) );
  OR2XLTH U895 ( .A(n722), .B(n795), .Y(n1072) );
  NAND2BXLTH U896 ( .AN(n1123), .B(n1102), .Y(n722) );
  NAND2XLTH U897 ( .A(n1149), .B(n1165), .Y(n907) );
  ADDFX1TH U898 ( .A(n572), .B(n603), .CI(n588), .CO(n444), .S(n445) );
  NOR2BXLTH U899 ( .AN(n1124), .B(n795), .Y(n572) );
  OAI22XLTH U900 ( .A0(n737), .A1(n1050), .B0(n736), .B1(n796), .Y(n588) );
  XNOR2X1TH U901 ( .A(n1113), .B(n1100), .Y(n749) );
  XNOR2X1TH U903 ( .A(n1112), .B(n1107), .Y(n631) );
  ADDFHXLTH U904 ( .A(n319), .B(n573), .CI(n462), .CO(n303), .S(n304) );
  NOR2BXLTH U905 ( .AN(n1110), .B(n1156), .Y(n462) );
  ADDFXLTH U906 ( .A(n555), .B(n289), .CI(n461), .CO(n275), .S(n276) );
  NOR2BXLTH U907 ( .AN(n1112), .B(n1156), .Y(n461) );
  ADDHX1TH U908 ( .A(n452), .B(n585), .CO(n434), .S(n435) );
  ADDFHXLTH U909 ( .A(n300), .B(n313), .CI(n557), .CO(n295), .S(n296) );
  ADDFHXLTH U910 ( .A(n317), .B(n315), .CI(n302), .CO(n297), .S(n298) );
  ADDFHXLTH U911 ( .A(n475), .B(n523), .CI(n287), .CO(n271), .S(n272) );
  OAI22XLTH U912 ( .A0(n629), .A1(n790), .B0(n630), .B1(n1048), .Y(n475) );
  NAND2XLTH U913 ( .A(n1110), .B(n1103), .Y(n916) );
  OR2XLTH U914 ( .A(n746), .B(n788), .Y(n886) );
  ADDFHXLTH U915 ( .A(n473), .B(n489), .CI(n252), .CO(n249), .S(n250) );
  OAI22XLTH U916 ( .A0(n627), .A1(n790), .B0(n628), .B1(n1048), .Y(n473) );
  ADDFHXLTH U917 ( .A(n598), .B(n423), .CI(n428), .CO(n418), .S(n419) );
  NAND2XLTH U918 ( .A(n425), .B(n430), .Y(n156) );
  NOR2XLTH U919 ( .A(n743), .B(n1099), .Y(n900) );
  CLKBUFX12TH U920 ( .A(a[13]), .Y(n1120) );
  NAND2XLTH U921 ( .A(n1119), .B(n1102), .Y(n935) );
  INVX5TH U922 ( .A(n96), .Y(n1129) );
  OR2XLTH U923 ( .A(n243), .B(n234), .Y(n923) );
  NAND2XLTH U924 ( .A(n243), .B(n234), .Y(n92) );
  OR2X1TH U925 ( .A(n278), .B(n291), .Y(n868) );
  NAND2XLTH U926 ( .A(n1112), .B(n1104), .Y(n891) );
  NAND2XLTH U927 ( .A(n1149), .B(n1159), .Y(n892) );
  XNOR2X1TH U928 ( .A(n1116), .B(n1102), .Y(n712) );
  NAND2XLTH U929 ( .A(n1120), .B(n1100), .Y(n963) );
  NAND2X1TH U930 ( .A(n1143), .B(n1165), .Y(n964) );
  INVX1TH U931 ( .A(n1120), .Y(n1143) );
  NAND2XLTH U932 ( .A(n1119), .B(n1101), .Y(n975) );
  XNOR2X1TH U933 ( .A(n1109), .B(n1106), .Y(n651) );
  NAND2XLTH U934 ( .A(n1137), .B(n71), .Y(n52) );
  NAND2XLTH U935 ( .A(n1032), .B(n1033), .Y(product_30_) );
  NAND2XLTH U936 ( .A(n69), .B(n51), .Y(n1032) );
  ADDFX2TH U937 ( .A(n592), .B(n357), .CI(n368), .CO(n352), .S(n353) );
  XNOR2X4TH U938 ( .A(n77), .B(n53), .Y(product_28_) );
  XNOR2X1TH U939 ( .A(n85), .B(n55), .Y(product_26_) );
  XNOR2X1TH U940 ( .A(n125), .B(n65), .Y(product_16_) );
  NAND2X4TH U941 ( .A(n778), .B(n795), .Y(n1051) );
  NAND2X4TH U942 ( .A(n775), .B(n792), .Y(n1052) );
  NAND2X4TH U943 ( .A(n777), .B(n794), .Y(n1053) );
  NAND2X4TH U944 ( .A(n776), .B(n793), .Y(n1054) );
  AND2XLTH U945 ( .A(n913), .B(n914), .Y(n1055) );
  NAND2XL U946 ( .A(n1117), .B(n1100), .Y(n949) );
  XNOR2XL U947 ( .A(n93), .B(n57), .Y(product_24_) );
  NAND2X5 U948 ( .A(n77), .B(n925), .Y(n1085) );
  NAND2X5 U949 ( .A(n985), .B(n79), .Y(n77) );
  NOR2X8 U950 ( .A(n1078), .B(n1077), .Y(n88) );
  NOR2X6 U951 ( .A(n1079), .B(n134), .Y(n970) );
  OAI22X1TH U952 ( .A0(n718), .A1(n795), .B0(n719), .B1(n1051), .Y(n569) );
  ADDFX2 U953 ( .A(n593), .B(n546), .CI(n875), .CO(n370), .S(n371) );
  CLKNAND2X4 U954 ( .A(n932), .B(n933), .Y(n746) );
  CLKNAND2X2 U955 ( .A(n339), .B(n352), .Y(n952) );
  CLKNAND2X2 U957 ( .A(n352), .B(n341), .Y(n954) );
  CLKNAND2X2 U958 ( .A(n339), .B(n341), .Y(n953) );
  CLKNAND2X2 U959 ( .A(n1110), .B(n1102), .Y(n1028) );
  CLKNAND2X2 U960 ( .A(n1152), .B(n1164), .Y(n1029) );
  CLKNAND2X2 U961 ( .A(n1146), .B(n1165), .Y(n961) );
  ADDFHX2TH U962 ( .A(n282), .B(n293), .CI(n280), .CO(n277), .S(n278) );
  CLKNAND2X4TH U963 ( .A(n278), .B(n291), .Y(n108) );
  INVX2TH U964 ( .A(n1123), .Y(n1069) );
  OR2XLTH U965 ( .A(n739), .B(n796), .Y(n1059) );
  NAND2BXLTH U966 ( .AN(n1123), .B(n1101), .Y(n739) );
  OAI22X1TH U967 ( .A0(n1090), .A1(n1050), .B0(n737), .B1(n796), .Y(n589) );
  NAND2X3TH U968 ( .A(n1063), .B(n1064), .Y(n602) );
  XNOR2XLTH U969 ( .A(n1123), .B(n1102), .Y(n721) );
  NOR2XLTH U970 ( .A(n704), .B(n1053), .Y(n1022) );
  CLKNAND2X2TH U971 ( .A(n1020), .B(n1021), .Y(n719) );
  ADDFHXLTH U972 ( .A(n509), .B(n477), .CI(n304), .CO(n301), .S(n302) );
  OAI22XLTH U973 ( .A0(n661), .A1(n792), .B0(n662), .B1(n1052), .Y(n509) );
  INVXLTH U974 ( .A(n1110), .Y(n1152) );
  OA21X2TH U975 ( .A0(n168), .A1(n166), .B0(n167), .Y(n1001) );
  NOR2X2TH U976 ( .A(n918), .B(n874), .Y(n168) );
  CLKNAND2X2TH U977 ( .A(n912), .B(n1055), .Y(n436) );
  OR2XLTH U978 ( .A(n1022), .B(n1023), .Y(n553) );
  OAI22XLTH U979 ( .A0(n748), .A1(n1099), .B0(n749), .B1(n788), .Y(n600) );
  NAND2XLTH U980 ( .A(n1108), .B(n1103), .Y(n909) );
  OAI22XLTH U981 ( .A0(n733), .A1(n796), .B0(n734), .B1(n1050), .Y(n585) );
  NAND2BXLTH U982 ( .AN(n1123), .B(n1103), .Y(n705) );
  ADDFHXLTH U983 ( .A(n541), .B(n493), .CI(n525), .CO(n299), .S(n300) );
  OAI22XLTH U984 ( .A0(n676), .A1(n793), .B0(n677), .B1(n1054), .Y(n525) );
  OAI22XLTH U985 ( .A0(n646), .A1(n791), .B0(n647), .B1(n1049), .Y(n493) );
  ADDFHXLTH U986 ( .A(n492), .B(n524), .CI(n303), .CO(n285), .S(n286) );
  ADDFHXLTH U987 ( .A(n491), .B(n507), .CI(n276), .CO(n273), .S(n274) );
  OAI22XLTH U988 ( .A0(n644), .A1(n791), .B0(n645), .B1(n1049), .Y(n491) );
  ADDFHXLTH U989 ( .A(n1130), .B(n490), .CI(n522), .CO(n261), .S(n262) );
  OAI22XLTH U990 ( .A0(n644), .A1(n1049), .B0(n643), .B1(n791), .Y(n490) );
  INVXLTH U991 ( .A(n263), .Y(n1130) );
  ADDFHXLTH U992 ( .A(n474), .B(n506), .CI(n275), .CO(n259), .S(n260) );
  ADDFHXLTH U993 ( .A(n536), .B(n568), .CI(n599), .CO(n428), .S(n429) );
  NOR2BXLTH U994 ( .AN(n1124), .B(n793), .Y(n536) );
  OAI22XLTH U995 ( .A0(n718), .A1(n1051), .B0(n717), .B1(n795), .Y(n568) );
  OR2XLTH U996 ( .A(n745), .B(n1099), .Y(n887) );
  INVX1TH U997 ( .A(n1109), .Y(n1153) );
  ADDFHXLTH U998 ( .A(n299), .B(n286), .CI(n556), .CO(n281), .S(n282) );
  OAI22XLTH U999 ( .A0(n706), .A1(n1051), .B0(n795), .B1(n1164), .Y(n556) );
  ADDFHXLTH U1000 ( .A(n285), .B(n274), .CI(n539), .CO(n269), .S(n270) );
  OAI22XLTH U1001 ( .A0(n689), .A1(n794), .B0(n690), .B1(n1053), .Y(n539) );
  ADDFHXLTH U1002 ( .A(n538), .B(n271), .CI(n258), .CO(n255), .S(n256) );
  ADDFHXLTH U1003 ( .A(n505), .B(n261), .CI(n259), .CO(n247), .S(n248) );
  OAI22XLTH U1004 ( .A0(n657), .A1(n792), .B0(n658), .B1(n1052), .Y(n505) );
  ADDFXLTH U1005 ( .A(n537), .B(n263), .CI(n460), .CO(n251), .S(n252) );
  NOR2BXLTH U1006 ( .AN(n1114), .B(n1156), .Y(n460) );
  ADDFHXLTH U1007 ( .A(n250), .B(n521), .CI(n248), .CO(n245), .S(n246) );
  OAI22XLTH U1008 ( .A0(n672), .A1(n793), .B0(n673), .B1(n1054), .Y(n521) );
  OAI22X1TH U1009 ( .A0(n716), .A1(n795), .B0(n717), .B1(n1051), .Y(n567) );
  OAI22X1TH U1010 ( .A0(n688), .A1(n793), .B0(n1054), .B1(n1159), .Y(n451) );
  NAND2BXLTH U1011 ( .AN(n1124), .B(n1104), .Y(n688) );
  ADDFHXLTH U1012 ( .A(n551), .B(n583), .CI(n535), .CO(n420), .S(n421) );
  OAI22XLTH U1014 ( .A0(n701), .A1(n794), .B0(n702), .B1(n1053), .Y(n551) );
  ADDFHXLTH U1015 ( .A(n518), .B(n550), .CI(n597), .CO(n414), .S(n415) );
  NOR2BXLTH U1016 ( .AN(n1124), .B(n792), .Y(n518) );
  NAND2XLTH U1017 ( .A(n886), .B(n887), .Y(n597) );
  NAND2XLTH U1018 ( .A(n1044), .B(n1045), .Y(n550) );
  ADDFHXLTH U1019 ( .A(n534), .B(n582), .CI(n566), .CO(n412), .S(n413) );
  OAI22XLTH U1020 ( .A0(n716), .A1(n1051), .B0(n715), .B1(n795), .Y(n566) );
  XNOR2X1TH U1021 ( .A(n1115), .B(n1101), .Y(n730) );
  ADDHXLTH U1022 ( .A(n450), .B(n596), .CO(n406), .S(n407) );
  OAI22XLTH U1023 ( .A0(n744), .A1(n1099), .B0(n745), .B1(n788), .Y(n596) );
  NAND2XLTH U1024 ( .A(n888), .B(n889), .Y(n450) );
  ADDFHXLTH U1025 ( .A(n526), .B(n494), .CI(n542), .CO(n315), .S(n316) );
  ADDFHXLTH U1026 ( .A(n527), .B(n495), .CI(n543), .CO(n331), .S(n332) );
  OAI22XLTH U1027 ( .A0(n648), .A1(n791), .B0(n649), .B1(n1049), .Y(n495) );
  OAI22XLTH U1028 ( .A0(n678), .A1(n793), .B0(n679), .B1(n1054), .Y(n527) );
  ADDFHXLTH U1029 ( .A(n270), .B(n279), .CI(n268), .CO(n265), .S(n266) );
  NAND2XLTH U1030 ( .A(n205), .B(n202), .Y(n71) );
  NAND2XLTH U1031 ( .A(n409), .B(n416), .Y(n148) );
  OAI22XLTH U1032 ( .A0(n714), .A1(n1051), .B0(n713), .B1(n795), .Y(n564) );
  ADDFHXLTH U1033 ( .A(n500), .B(n532), .CI(n580), .CO(n396), .S(n397) );
  NOR2BXLTH U1034 ( .AN(n1124), .B(n791), .Y(n500) );
  NAND2XLTH U1035 ( .A(n1040), .B(n1041), .Y(n580) );
  XNOR2X1TH U1036 ( .A(n1117), .B(n1102), .Y(n711) );
  XNOR2X1TH U1037 ( .A(n1108), .B(n1107), .Y(n635) );
  ADDFHXLTH U1038 ( .A(n510), .B(n558), .CI(n333), .CO(n313), .S(n314) );
  OAI22XLTH U1039 ( .A0(n663), .A1(n1052), .B0(n662), .B1(n792), .Y(n510) );
  ADDFHXLTH U1040 ( .A(n511), .B(n559), .CI(n334), .CO(n329), .S(n330) );
  OAI22XLTH U1042 ( .A0(n663), .A1(n792), .B0(n664), .B1(n1052), .Y(n511) );
  ADDFHXLTH U1043 ( .A(n348), .B(n346), .CI(n332), .CO(n327), .S(n328) );
  OAI22XLTH U1044 ( .A0(n727), .A1(n1050), .B0(n726), .B1(n796), .Y(n578) );
  CLKAND2X4TH U1045 ( .A(n1086), .B(n84), .Y(n80) );
  OR2XLTH U1046 ( .A(n265), .B(n254), .Y(n876) );
  NAND2XLTH U1047 ( .A(n265), .B(n254), .Y(n100) );
  AND2X6 U1048 ( .A(n93), .B(n923), .Y(n1078) );
  OAI22XLTH U1049 ( .A0(n712), .A1(n795), .B0(n713), .B1(n1051), .Y(n563) );
  ADDFHXLTH U1050 ( .A(n497), .B(n577), .CI(n529), .CO(n358), .S(n359) );
  ADDFHXLTH U1051 ( .A(n327), .B(n312), .CI(n325), .CO(n307), .S(n308) );
  ADDFX1TH U1052 ( .A(n349), .B(n358), .CI(n347), .CO(n342), .S(n343) );
  XOR2X1TH U1053 ( .A(n96), .B(n58), .Y(product_23_) );
  NAND2XLTH U1054 ( .A(n1126), .B(n1139), .Y(n1033) );
  INVXLTH U1055 ( .A(n51), .Y(n1139) );
  NOR2XLTH U1056 ( .A(n389), .B(n398), .Y(n139) );
  NAND2XLTH U1057 ( .A(n353), .B(n355), .Y(n939) );
  NAND2XLTH U1058 ( .A(n366), .B(n355), .Y(n940) );
  NAND2XLTH U1059 ( .A(n353), .B(n366), .Y(n938) );
  NAND2XLTH U1060 ( .A(n1131), .B(n127), .Y(n66) );
  NAND2XLTH U1061 ( .A(n1132), .B(n119), .Y(n64) );
  AND2XLTH U1063 ( .A(n1121), .B(n1101), .Y(n1057) );
  NAND2XLTH U1064 ( .A(n879), .B(n880), .Y(product_19_) );
  INVXLTH U1066 ( .A(n70), .Y(n1137) );
  NAND2XLTH U1067 ( .A(n924), .B(n84), .Y(n55) );
  OR2XLTH U1068 ( .A(n753), .B(n1099), .Y(n1066) );
  OAI22XLTH U1069 ( .A0(n746), .A1(n1099), .B0(n747), .B1(n788), .Y(n598) );
  OAI22XLTH U1070 ( .A0(n748), .A1(n788), .B0(n747), .B1(n1099), .Y(n599) );
  NOR2X8 U1071 ( .A(n1076), .B(n1075), .Y(n96) );
  AOI21BX4 U1072 ( .A0(n117), .A1(n863), .B0N(n116), .Y(n112) );
  NOR2X4 U1073 ( .A(n292), .B(n305), .Y(n110) );
  AOI21BX4 U1074 ( .A0(n125), .A1(n862), .B0N(n124), .Y(n120) );
  CLKNAND2X4 U1075 ( .A(n884), .B(n885), .Y(n747) );
  BUFX12 U1076 ( .A(a[3]), .Y(n1110) );
  NAND2X4 U1077 ( .A(n902), .B(n903), .Y(n716) );
  BUFX5 U1078 ( .A(n1056), .Y(n1124) );
  CLKNAND2X4TH U1079 ( .A(n1136), .B(n1165), .Y(n950) );
  CLKNAND2X4TH U1080 ( .A(n351), .B(n364), .Y(n127) );
  NOR2X4TH U1081 ( .A(n277), .B(n266), .Y(n102) );
  CLKNAND2X2 U1082 ( .A(n277), .B(n266), .Y(n103) );
  OR2XLTH U1083 ( .A(n1050), .B(n1160), .Y(n1060) );
  CLKNAND2X4TH U1084 ( .A(n1067), .B(n1068), .Y(n586) );
  CLKNAND2X2 U1085 ( .A(n1118), .B(n1100), .Y(n960) );
  ADDFHXLTH U1086 ( .A(n1161), .B(n464), .CI(n479), .CO(n333), .S(n334) );
  CLKNAND2X2 U1087 ( .A(n1144), .B(n1160), .Y(n976) );
  CLKNAND2X2 U1088 ( .A(n112), .B(n1133), .Y(n879) );
  NAND2X1 U1089 ( .A(n1014), .B(n87), .Y(n56) );
  CLKNAND2X2 U1090 ( .A(n365), .B(n376), .Y(n132) );
  NOR2X4TH U1091 ( .A(n970), .B(n927), .Y(n996) );
  NOR2X4 U1092 ( .A(n351), .B(n364), .Y(n126) );
  NAND2XLTH U1093 ( .A(n1123), .B(n1100), .Y(n1070) );
  NAND2XLTH U1094 ( .A(n1069), .B(n1165), .Y(n1071) );
  NAND2BXLTH U1095 ( .AN(n1123), .B(n1100), .Y(n756) );
  OR2XLTH U1096 ( .A(n753), .B(n788), .Y(n1062) );
  OR2XLTH U1097 ( .A(n752), .B(n1099), .Y(n1061) );
  NAND2XLTH U1098 ( .A(n605), .B(n590), .Y(n180) );
  OR2XLTH U1099 ( .A(n751), .B(n788), .Y(n1064) );
  XNOR2X1TH U1100 ( .A(n1110), .B(n1101), .Y(n735) );
  NAND2XLTH U1101 ( .A(n1112), .B(n1100), .Y(n906) );
  NAND2XLTH U1102 ( .A(n1109), .B(n1102), .Y(n1020) );
  XNOR2X1TH U1103 ( .A(n1114), .B(n1106), .Y(n646) );
  XNOR2X1TH U1104 ( .A(n1115), .B(n1106), .Y(n645) );
  XNOR2X1TH U1105 ( .A(n1116), .B(n1106), .Y(n644) );
  XNOR2X1TH U1106 ( .A(n1119), .B(n1104), .Y(n675) );
  XNOR2X1TH U1107 ( .A(n1120), .B(n1104), .Y(n674) );
  XNOR2X1TH U1108 ( .A(n1114), .B(n1100), .Y(n748) );
  NAND2XLTH U1109 ( .A(n441), .B(n444), .Y(n167) );
  NOR2XLTH U1110 ( .A(n441), .B(n444), .Y(n166) );
  XNOR2X1TH U1111 ( .A(n1119), .B(n1105), .Y(n658) );
  XNOR2X1TH U1112 ( .A(n1117), .B(n1106), .Y(n643) );
  XNOR2X1TH U1113 ( .A(n1120), .B(n1105), .Y(n657) );
  XNOR2X1TH U1114 ( .A(n1117), .B(n1107), .Y(n626) );
  XNOR2X1TH U1115 ( .A(n1120), .B(n1106), .Y(n640) );
  ADDFHXLTH U1116 ( .A(n476), .B(n288), .CI(n301), .CO(n283), .S(n284) );
  CLKINVX2TH U1117 ( .A(n1103), .Y(n1163) );
  XNOR2X1TH U1118 ( .A(n1119), .B(n1103), .Y(n692) );
  CLKINVX2TH U1119 ( .A(n1102), .Y(n1164) );
  INVXLTH U1120 ( .A(n319), .Y(n1161) );
  NAND2BXLTH U1121 ( .AN(n1115), .B(n1165), .Y(n885) );
  NAND2BXLTH U1122 ( .AN(n1116), .B(n1165), .Y(n933) );
  NOR2XLTH U1123 ( .A(n425), .B(n430), .Y(n155) );
  NAND2XLTH U1124 ( .A(n1114), .B(n1101), .Y(n897) );
  NAND2XLTH U1125 ( .A(n1148), .B(n1160), .Y(n898) );
  INVXLTH U1126 ( .A(n1114), .Y(n1148) );
  NAND2XLTH U1127 ( .A(n1112), .B(n1102), .Y(n902) );
  CLKNAND2X4TH U1128 ( .A(n1149), .B(n1164), .Y(n903) );
  NAND2BXLTH U1129 ( .AN(n1124), .B(n1105), .Y(n671) );
  CLKBUFX6TH U1130 ( .A(b[5]), .Y(n1102) );
  CLKBUFX6TH U1131 ( .A(b[7]), .Y(n1103) );
  XNOR2X1TH U1132 ( .A(n1119), .B(n1107), .Y(n624) );
  XNOR2X1TH U1133 ( .A(n1120), .B(n1107), .Y(n623) );
  ADDFXLTH U1134 ( .A(n501), .B(n223), .CI(n458), .CO(n215), .S(n216) );
  NOR2BXLTH U1135 ( .AN(n1118), .B(n1156), .Y(n458) );
  CLKINVX2TH U1136 ( .A(n1104), .Y(n1159) );
  XNOR2X1TH U1137 ( .A(n1119), .B(n1106), .Y(n641) );
  CLKBUFX6TH U1138 ( .A(b[9]), .Y(n1104) );
  CLKBUFX6TH U1139 ( .A(b[11]), .Y(n1105) );
  XNOR2X1TH U1140 ( .A(n1121), .B(n1105), .Y(n656) );
  ADDFHXLTH U1141 ( .A(n1147), .B(n472), .CI(n504), .CO(n239), .S(n240) );
  OAI22XLTH U1142 ( .A0(n627), .A1(n1048), .B0(n626), .B1(n790), .Y(n472) );
  INVXLTH U1143 ( .A(n241), .Y(n1147) );
  ADDFXLTH U1144 ( .A(n519), .B(n241), .CI(n459), .CO(n231), .S(n232) );
  NOR2BXLTH U1145 ( .AN(n1116), .B(n1156), .Y(n459) );
  ADDFHXLTH U1146 ( .A(n487), .B(n471), .CI(n232), .CO(n229), .S(n230) );
  OAI22XLTH U1147 ( .A0(n625), .A1(n790), .B0(n626), .B1(n1048), .Y(n471) );
  ADDFHXLTH U1148 ( .A(n1138), .B(n486), .CI(n470), .CO(n221), .S(n222) );
  INVXLTH U1149 ( .A(n223), .Y(n1138) );
  ADDFHXLTH U1150 ( .A(n311), .B(n298), .CI(n296), .CO(n293), .S(n294) );
  ADDFHXLTH U1151 ( .A(n262), .B(n273), .CI(n260), .CO(n257), .S(n258) );
  ADDFHXLTH U1152 ( .A(n297), .B(n284), .CI(n295), .CO(n279), .S(n280) );
  ADDFHXLTH U1153 ( .A(n272), .B(n283), .CI(n281), .CO(n267), .S(n268) );
  XNOR2X1TH U1154 ( .A(n1121), .B(n1107), .Y(n622) );
  ADDFHXLTH U1155 ( .A(n1161), .B(n463), .CI(n478), .CO(n317), .S(n318) );
  NOR2XLTH U1156 ( .A(n1153), .B(n1156), .Y(n463) );
  XNOR2X1TH U1157 ( .A(n1115), .B(n1105), .Y(n662) );
  XNOR2X1TH U1158 ( .A(n1109), .B(n1107), .Y(n634) );
  XNOR2X1TH U1159 ( .A(n1114), .B(n1105), .Y(n663) );
  CLKBUFX6TH U1160 ( .A(b[3]), .Y(n1101) );
  CLKBUFX6TH U1161 ( .A(b[15]), .Y(n1107) );
  INVX4TH U1162 ( .A(n1107), .Y(n1156) );
  CLKBUFX6TH U1163 ( .A(b[13]), .Y(n1106) );
  XOR2XLTH U1164 ( .A(b[14]), .B(n1107), .Y(n773) );
  CLKBUFX6TH U1165 ( .A(b[1]), .Y(n1100) );
  INVX4TH U1166 ( .A(n1097), .Y(n790) );
  XOR2XLTH U1167 ( .A(b[14]), .B(n1106), .Y(n1097) );
  INVX5TH U1168 ( .A(n1091), .Y(n795) );
  XOR2XLTH U1169 ( .A(b[4]), .B(n1101), .Y(n1091) );
  XOR2XLTH U1170 ( .A(b[4]), .B(n1102), .Y(n778) );
  XOR2XLTH U1171 ( .A(b[8]), .B(n1103), .Y(n1095) );
  XOR2XLTH U1172 ( .A(b[8]), .B(n1104), .Y(n776) );
  INVX5TH U1173 ( .A(n1092), .Y(n794) );
  XOR2XLTH U1174 ( .A(b[6]), .B(n1102), .Y(n1092) );
  XOR2XLTH U1175 ( .A(b[6]), .B(n1103), .Y(n777) );
  INVXLTH U1176 ( .A(n112), .Y(n1125) );
  INVXLTH U1177 ( .A(n110), .Y(n1134) );
  XOR2XLTH U1178 ( .A(b[12]), .B(n1105), .Y(n1096) );
  XOR2XLTH U1179 ( .A(b[12]), .B(n1106), .Y(n774) );
  ADDFHXLTH U1180 ( .A(n469), .B(n216), .CI(n221), .CO(n213), .S(n214) );
  OAI22XLTH U1181 ( .A0(n623), .A1(n790), .B0(n624), .B1(n1048), .Y(n469) );
  CLKINVX1TH U1182 ( .A(n1106), .Y(n1157) );
  ADDFHXLTH U1183 ( .A(n1145), .B(n468), .CI(n215), .CO(n207), .S(n208) );
  INVXLTH U1184 ( .A(n209), .Y(n1145) );
  OAI22XLTH U1185 ( .A0(n623), .A1(n1048), .B0(n622), .B1(n790), .Y(n468) );
  ADDFHXLTH U1186 ( .A(n249), .B(n520), .CI(n247), .CO(n235), .S(n236) );
  ADDFHXLTH U1187 ( .A(n488), .B(n251), .CI(n240), .CO(n237), .S(n238) );
  OAI22XLTH U1188 ( .A0(n642), .A1(n1049), .B0(n641), .B1(n791), .Y(n488) );
  CLKINVX1TH U1189 ( .A(n1105), .Y(n1158) );
  INVX5TH U1190 ( .A(n1094), .Y(n792) );
  XOR2XLTH U1191 ( .A(b[10]), .B(n1104), .Y(n1094) );
  XOR2XLTH U1192 ( .A(b[10]), .B(n1105), .Y(n775) );
  ADDFHXLTH U1193 ( .A(n239), .B(n230), .CI(n503), .CO(n227), .S(n228) );
  OAI22XLTH U1194 ( .A0(n655), .A1(n792), .B0(n656), .B1(n1052), .Y(n503) );
  ADDFHXLTH U1195 ( .A(n231), .B(n222), .CI(n229), .CO(n219), .S(n220) );
  ADDFHXLTH U1196 ( .A(n257), .B(n255), .CI(n246), .CO(n243), .S(n244) );
  ADDFHXLTH U1197 ( .A(n269), .B(n256), .CI(n267), .CO(n253), .S(n254) );
  ADDFHXLTH U1198 ( .A(n238), .B(n245), .CI(n236), .CO(n233), .S(n234) );
  NOR2XLTH U1199 ( .A(n1142), .B(n1156), .Y(n456) );
  ADDFXLTH U1200 ( .A(n483), .B(n209), .CI(n457), .CO(n203), .S(n204) );
  NOR2BXLTH U1201 ( .AN(n1120), .B(n1156), .Y(n457) );
  ADDFHXLTH U1202 ( .A(n204), .B(n207), .CI(n467), .CO(n201), .S(n202) );
  OAI22XLTH U1203 ( .A0(n621), .A1(n790), .B0(n622), .B1(n1048), .Y(n467) );
  NOR2XLTH U1204 ( .A(n205), .B(n202), .Y(n70) );
  INVX3TH U1205 ( .A(n1100), .Y(n1165) );
  ADDFHXLTH U1206 ( .A(n318), .B(n331), .CI(n316), .CO(n311), .S(n312) );
  CLKINVX2TH U1207 ( .A(n1101), .Y(n1160) );
  XOR2XLTH U1208 ( .A(b[2]), .B(n1101), .Y(n779) );
  INVX5TH U1209 ( .A(n1093), .Y(n796) );
  XOR2XLTH U1210 ( .A(b[2]), .B(n1100), .Y(n1093) );
  ADDFHXLTH U1211 ( .A(n528), .B(n512), .CI(n560), .CO(n346), .S(n347) );
  NAND2XLTH U1212 ( .A(n919), .B(n920), .Y(n560) );
  ADDFHXLTH U1213 ( .A(n465), .B(n496), .CI(n544), .CO(n348), .S(n349) );
  NOR2BXLTH U1214 ( .AN(n1124), .B(n1156), .Y(n465) );
  OAI22XLTH U1215 ( .A0(n650), .A1(n1049), .B0(n649), .B1(n791), .Y(n496) );
  ADDFHXLTH U1216 ( .A(n533), .B(n549), .CI(n517), .CO(n404), .S(n405) );
  OAI22XLTH U1217 ( .A0(n684), .A1(n793), .B0(n685), .B1(n1054), .Y(n533) );
  ADDFHXLTH U1218 ( .A(n581), .B(n565), .CI(n407), .CO(n402), .S(n403) );
  ADDFHXLTH U1219 ( .A(n564), .B(n595), .CI(n548), .CO(n394), .S(n395) );
  OR2XLTH U1220 ( .A(n899), .B(n900), .Y(n595) );
  INVXLTH U1221 ( .A(n579), .Y(n1140) );
  ADDFHXLTH U1222 ( .A(n545), .B(n561), .CI(n481), .CO(n360), .S(n361) );
  OAI22XLTH U1223 ( .A0(n695), .A1(n794), .B0(n696), .B1(n1053), .Y(n545) );
  OAI22XLTH U1224 ( .A0(n680), .A1(n793), .B0(n681), .B1(n1054), .Y(n529) );
  OAI22XLTH U1225 ( .A0(n650), .A1(n791), .B0(n651), .B1(n1049), .Y(n497) );
  BUFX4TH U1226 ( .A(n1162), .Y(n1099) );
  INVXLTH U1227 ( .A(b[0]), .Y(n1162) );
  INVX4TH U1228 ( .A(n1098), .Y(n788) );
  AND2XLTH U1229 ( .A(n780), .B(n1099), .Y(n1098) );
  XOR2XLTH U1230 ( .A(b[0]), .B(n1100), .Y(n780) );
  INVXLTH U1231 ( .A(n1122), .Y(n1141) );
  ADDFHXLTH U1232 ( .A(n516), .B(n406), .CI(n397), .CO(n392), .S(n393) );
  ADDFHXLTH U1233 ( .A(n515), .B(n547), .CI(n594), .CO(n382), .S(n383) );
  OAI22XLTH U1234 ( .A0(n697), .A1(n794), .B0(n698), .B1(n1053), .Y(n547) );
  NAND2XLTH U1235 ( .A(n1034), .B(n1035), .Y(n594) );
  OAI22XLTH U1236 ( .A0(n667), .A1(n792), .B0(n668), .B1(n1052), .Y(n515) );
  ADDFHXLTH U1237 ( .A(n482), .B(n514), .CI(n562), .CO(n374), .S(n375) );
  NOR2BXLTH U1238 ( .AN(n1124), .B(n790), .Y(n482) );
  ADDFHXLTH U1239 ( .A(n498), .B(n530), .CI(n578), .CO(n372), .S(n373) );
  OAI22XLTH U1240 ( .A0(n682), .A1(n1054), .B0(n681), .B1(n793), .Y(n530) );
  ADDFHXLTH U1241 ( .A(n563), .B(n531), .CI(n499), .CO(n384), .S(n385) );
  OAI22XLTH U1242 ( .A0(n682), .A1(n793), .B0(n683), .B1(n1054), .Y(n531) );
  AND2XLTH U1243 ( .A(n1047), .B(n579), .Y(n875) );
  ADDFHXLTH U1244 ( .A(n485), .B(n214), .CI(n219), .CO(n211), .S(n212) );
  OAI22XLTH U1245 ( .A0(n638), .A1(n791), .B0(n639), .B1(n1049), .Y(n485) );
  ADDFHXLTH U1246 ( .A(n208), .B(n484), .CI(n213), .CO(n205), .S(n206) );
  ADDFHXLTH U1247 ( .A(n237), .B(n228), .CI(n235), .CO(n225), .S(n226) );
  ADDFHXLTH U1248 ( .A(n502), .B(n220), .CI(n227), .CO(n217), .S(n218) );
  OR2XLTH U1249 ( .A(n253), .B(n244), .Y(n867) );
  NAND2X1TH U1250 ( .A(n253), .B(n244), .Y(n95) );
  OR2XLTH U1251 ( .A(n217), .B(n212), .Y(n1058) );
  NAND2XLTH U1252 ( .A(n217), .B(n212), .Y(n79) );
  INVXLTH U1253 ( .A(n92), .Y(n1077) );
  OR2XLTH U1254 ( .A(n233), .B(n226), .Y(n1014) );
  NAND2X1TH U1255 ( .A(n233), .B(n226), .Y(n87) );
  NAND2XLTH U1256 ( .A(n923), .B(n92), .Y(n57) );
  NAND2BXLTH U1257 ( .AN(n1012), .B(n68), .Y(n51) );
  NAND2XLTH U1258 ( .A(n199), .B(n201), .Y(n68) );
  NOR2XLTH U1259 ( .A(n199), .B(n201), .Y(n1012) );
  XNOR3XLTH U1260 ( .A(n456), .B(n203), .C(n994), .Y(n199) );
  ADDFHXLTH U1262 ( .A(n329), .B(n314), .CI(n574), .CO(n309), .S(n310) );
  ADDFHXLTH U1263 ( .A(n344), .B(n575), .CI(n330), .CO(n325), .S(n326) );
  ADDFHXLTH U1264 ( .A(n342), .B(n328), .CI(n340), .CO(n323), .S(n324) );
  ADDFX1TH U1265 ( .A(n363), .B(n374), .CI(n372), .CO(n356), .S(n357) );
  NAND2XLTH U1266 ( .A(n1017), .B(n1018), .Y(n387) );
  NAND2XLTH U1267 ( .A(n1155), .B(n579), .Y(n1018) );
  ADDFHXLTH U1268 ( .A(n383), .B(n385), .CI(n392), .CO(n378), .S(n379) );
  ADDFHXLTH U1269 ( .A(n375), .B(n382), .CI(n373), .CO(n368), .S(n369) );
  ADDFX1TH U1270 ( .A(n384), .B(n371), .CI(n380), .CO(n366), .S(n367) );
  INVX1TH U1271 ( .A(n80), .Y(n1127) );
  OR2XLTH U1272 ( .A(n211), .B(n206), .Y(n925) );
  NAND2XLTH U1274 ( .A(n211), .B(n206), .Y(n76) );
  OR2XLTH U1275 ( .A(n225), .B(n218), .Y(n924) );
  NAND2XLTH U1276 ( .A(n225), .B(n218), .Y(n84) );
  NAND2XLTH U1277 ( .A(n1135), .B(n103), .Y(n60) );
  NAND2XLTH U1278 ( .A(n867), .B(n95), .Y(n58) );
  NAND2XLTH U1279 ( .A(n1058), .B(n79), .Y(n54) );
  NAND2XLTH U1280 ( .A(n343), .B(n354), .Y(n1037) );
  NAND2XLTH U1281 ( .A(n343), .B(n356), .Y(n1038) );
  NAND2XLTH U1282 ( .A(n389), .B(n398), .Y(n140) );
  CLKXOR2X2TH U1283 ( .A(n937), .B(n353), .Y(n351) );
  XOR2X2TH U1284 ( .A(n355), .B(n366), .Y(n937) );
  ADDFX1TH U1285 ( .A(n369), .B(n378), .CI(n367), .CO(n364), .S(n365) );
  NAND2XLTH U1286 ( .A(n925), .B(n76), .Y(n53) );
  OR2XLTH U1287 ( .A(n306), .B(n321), .Y(n863) );
  INVXLTH U1288 ( .A(n126), .Y(n1131) );
  OAI22XLTH U1289 ( .A0(n636), .A1(n1048), .B0(n635), .B1(n790), .Y(n481) );
  OAI22XLTH U1290 ( .A0(n635), .A1(n1048), .B0(n634), .B1(n790), .Y(n480) );
  OAI22XLTH U1291 ( .A0(n631), .A1(n1048), .B0(n630), .B1(n790), .Y(n476) );
  OAI22XLTH U1292 ( .A0(n629), .A1(n1048), .B0(n628), .B1(n790), .Y(n474) );
  OAI22XLTH U1293 ( .A0(n625), .A1(n1048), .B0(n624), .B1(n790), .Y(n470) );
  OAI22XLTH U1294 ( .A0(n689), .A1(n1053), .B0(n794), .B1(n1163), .Y(n538) );
  OAI22XLTH U1295 ( .A0(n699), .A1(n1053), .B0(n698), .B1(n794), .Y(n548) );
  OAI22XLTH U1296 ( .A0(n697), .A1(n1053), .B0(n696), .B1(n794), .Y(n546) );
  OAI22XLTH U1297 ( .A0(n703), .A1(n1053), .B0(n702), .B1(n794), .Y(n552) );
  OAI22XLTH U1298 ( .A0(n705), .A1(n794), .B0(n1053), .B1(n1163), .Y(n452) );
  OAI22XLTH U1299 ( .A0(n655), .A1(n1052), .B0(n792), .B1(n1158), .Y(n502) );
  OAI22XLTH U1300 ( .A0(n667), .A1(n1052), .B0(n666), .B1(n792), .Y(n514) );
  OAI22XLTH U1301 ( .A0(n665), .A1(n1052), .B0(n664), .B1(n792), .Y(n512) );
  OAI22XLTH U1302 ( .A0(n669), .A1(n1052), .B0(n668), .B1(n792), .Y(n516) );
  OAI22XLTH U1303 ( .A0(n670), .A1(n1052), .B0(n669), .B1(n792), .Y(n517) );
  OAI22XLTH U1304 ( .A0(n672), .A1(n1054), .B0(n793), .B1(n1159), .Y(n520) );
  OAI22XLTH U1305 ( .A0(n687), .A1(n1054), .B0(n686), .B1(n793), .Y(n535) );
  OAI22XLTH U1306 ( .A0(n680), .A1(n1054), .B0(n679), .B1(n793), .Y(n528) );
  OAI22XLTH U1307 ( .A0(n678), .A1(n1054), .B0(n677), .B1(n793), .Y(n526) );
  OAI22XLTH U1308 ( .A0(n686), .A1(n1054), .B0(n685), .B1(n793), .Y(n534) );
  INVX5TH U1309 ( .A(n1095), .Y(n793) );
  OAI22XLTH U1310 ( .A0(n638), .A1(n1049), .B0(n791), .B1(n1157), .Y(n484) );
  OAI22XLTH U1311 ( .A0(n652), .A1(n1049), .B0(n651), .B1(n791), .Y(n498) );
  OAI22XLTH U1312 ( .A0(n653), .A1(n1049), .B0(n652), .B1(n791), .Y(n499) );
  OAI22XLTH U1313 ( .A0(n648), .A1(n1049), .B0(n647), .B1(n791), .Y(n494) );
  OAI22XLTH U1314 ( .A0(n646), .A1(n1049), .B0(n645), .B1(n791), .Y(n492) );
  INVX5TH U1315 ( .A(n1096), .Y(n791) );
  OAI22X1 U1316 ( .A0(n720), .A1(n1051), .B0(n719), .B1(n795), .Y(n570) );
  XOR2X4 U1317 ( .A(n453), .B(n602), .Y(n443) );
  NAND2XLTH U1318 ( .A(n439), .B(n873), .Y(n913) );
  OR2X4 U1319 ( .A(n431), .B(n436), .Y(n1088) );
  OR2XLTH U1320 ( .A(n735), .B(n1050), .Y(n1067) );
  OR2XLTH U1321 ( .A(n734), .B(n796), .Y(n1068) );
  ADDFHX4 U1322 ( .A(n554), .B(n586), .CI(n570), .CO(n438), .S(n439) );
  OR2XLTH U1323 ( .A(n1051), .B(n1164), .Y(n1073) );
  BUFX10 U1324 ( .A(a[6]), .Y(n1113) );
  AND2X6 U1325 ( .A(n1085), .B(n76), .Y(n72) );
  NOR2X4 U1326 ( .A(n941), .B(n926), .Y(n998) );
  AND2XLTH U1327 ( .A(n399), .B(n408), .Y(n926) );
  ADDFHX2 U1328 ( .A(n587), .B(n571), .CI(n443), .CO(n440), .S(n441) );
  NAND2XLTH U1329 ( .A(n1116), .B(n1100), .Y(n932) );
  XNOR2X1TH U1330 ( .A(n1114), .B(n1107), .Y(n629) );
  NAND2XLTH U1331 ( .A(n876), .B(n100), .Y(n59) );
  BUFX8 U1332 ( .A(a[7]), .Y(n1114) );
  NAND2X1TH U1333 ( .A(n292), .B(n305), .Y(n111) );
  XNOR2X1TH U1334 ( .A(n1111), .B(n1102), .Y(n717) );
  NAND2XLTH U1335 ( .A(n1115), .B(n1100), .Y(n884) );
  XNOR2X1TH U1336 ( .A(n1115), .B(n1107), .Y(n628) );
  XNOR2X1TH U1337 ( .A(n1116), .B(n1107), .Y(n627) );
  XNOR2X1TH U1338 ( .A(n1121), .B(n1106), .Y(n639) );
  INVXLTH U1339 ( .A(n100), .Y(n1075) );
  NOR2BXLTH U1340 ( .AN(n1113), .B(n1156), .Y(n263) );
  XNOR2X1 U1341 ( .A(n1114), .B(n1102), .Y(n714) );
  INVXLTH U1342 ( .A(n1117), .Y(n1136) );
  AND2XLTH U1343 ( .A(n1142), .B(n1160), .Y(n1081) );
  NAND2XLTH U1344 ( .A(n862), .B(n124), .Y(n65) );
  NAND2XLTH U1345 ( .A(n868), .B(n108), .Y(n61) );
  INVXLTH U1346 ( .A(n102), .Y(n1135) );
  OA21X4 U1347 ( .A0(n998), .A1(n139), .B0(n140), .Y(n1079) );
  OA21X4 U1348 ( .A0(n996), .A1(n131), .B0(n132), .Y(n128) );
  AND2XLTH U1349 ( .A(n377), .B(n388), .Y(n927) );
  OA21X4 U1350 ( .A0(n999), .A1(n155), .B0(n156), .Y(n152) );
  NAND2XLTH U1351 ( .A(n354), .B(n356), .Y(n1039) );
  OA21X4 U1352 ( .A0(n176), .A1(n174), .B0(n175), .Y(n1080) );
  AND2XLTH U1353 ( .A(n451), .B(n567), .Y(n1013) );
  OAI22XLTH U1354 ( .A0(n684), .A1(n1054), .B0(n683), .B1(n793), .Y(n532) );
  OAI22XLTH U1355 ( .A0(n695), .A1(n1053), .B0(n694), .B1(n794), .Y(n544) );
  NOR2XLTH U1356 ( .A(n744), .B(n788), .Y(n899) );
  OAI22XLTH U1357 ( .A0(n699), .A1(n794), .B0(n700), .B1(n1053), .Y(n549) );
  OAI22XLTH U1358 ( .A0(n714), .A1(n795), .B0(n715), .B1(n1051), .Y(n565) );
  OAI22XLTH U1359 ( .A0(n631), .A1(n790), .B0(n632), .B1(n1048), .Y(n477) );
  OAI22XLTH U1360 ( .A0(n693), .A1(n1053), .B0(n692), .B1(n794), .Y(n542) );
  OAI22XLTH U1361 ( .A0(n693), .A1(n794), .B0(n694), .B1(n1053), .Y(n543) );
  OAI22XLTH U1362 ( .A0(n633), .A1(n1048), .B0(n632), .B1(n790), .Y(n478) );
  OAI22XLTH U1363 ( .A0(n674), .A1(n1054), .B0(n673), .B1(n793), .Y(n522) );
  OAI22XLTH U1364 ( .A0(n676), .A1(n1054), .B0(n675), .B1(n793), .Y(n524) );
  OAI22XLTH U1365 ( .A0(n659), .A1(n1052), .B0(n658), .B1(n792), .Y(n506) );
  NOR2BXLTH U1366 ( .AN(n1111), .B(n1156), .Y(n289) );
  OAI22XLTH U1367 ( .A0(n659), .A1(n792), .B0(n660), .B1(n1052), .Y(n507) );
  OAI22XLTH U1368 ( .A0(n674), .A1(n793), .B0(n675), .B1(n1054), .Y(n523) );
  OAI22XLTH U1369 ( .A0(n640), .A1(n791), .B0(n641), .B1(n1049), .Y(n487) );
  NOR2BXLTH U1370 ( .AN(n1115), .B(n1156), .Y(n241) );
  OAI22XLTH U1371 ( .A0(n657), .A1(n1052), .B0(n656), .B1(n792), .Y(n504) );
  OAI22XLTH U1372 ( .A0(n642), .A1(n791), .B0(n643), .B1(n1049), .Y(n489) );
  OAI22XLTH U1373 ( .A0(n640), .A1(n1049), .B0(n639), .B1(n791), .Y(n486) );
  NOR2BXLTH U1374 ( .AN(n1117), .B(n1156), .Y(n223) );
  NOR2BXLTH U1375 ( .AN(n1119), .B(n1156), .Y(n209) );
  OAI22XLTH U1376 ( .A0(n621), .A1(n1048), .B0(n790), .B1(n1156), .Y(n994) );
  XNOR2X1TH U1377 ( .A(n1113), .B(n1101), .Y(n732) );
  XNOR2X1TH U1378 ( .A(n1109), .B(n1101), .Y(n736) );
  XNOR2X1TH U1379 ( .A(n1109), .B(n1103), .Y(n702) );
  XNOR2X1TH U1380 ( .A(n1112), .B(n1101), .Y(n733) );
  XNOR2X1TH U1381 ( .A(n1111), .B(n1103), .Y(n700) );
  XNOR2XLTH U1382 ( .A(n1123), .B(n1101), .Y(n1090) );
  XNOR2XLTH U1383 ( .A(n1123), .B(n1103), .Y(n704) );
  NAND2BX1TH U1384 ( .AN(n1124), .B(n1106), .Y(n654) );
  XNOR2X1TH U1385 ( .A(n1108), .B(n1105), .Y(n669) );
  XNOR2X1TH U1386 ( .A(n1113), .B(n1102), .Y(n715) );
  XNOR2X1TH U1387 ( .A(n1113), .B(n1103), .Y(n698) );
  XNOR2X1TH U1388 ( .A(n1113), .B(n1104), .Y(n681) );
  XNOR2X1TH U1389 ( .A(n1113), .B(n1105), .Y(n664) );
  XNOR2X1TH U1390 ( .A(n1112), .B(n1103), .Y(n699) );
  XNOR2X1TH U1391 ( .A(n1110), .B(n1104), .Y(n684) );
  XNOR2X1TH U1392 ( .A(n1116), .B(n1103), .Y(n695) );
  XNOR2X1TH U1393 ( .A(n1114), .B(n1103), .Y(n697) );
  XNOR2X1TH U1394 ( .A(n1114), .B(n1104), .Y(n680) );
  XNOR2X1TH U1395 ( .A(n1110), .B(n1105), .Y(n667) );
  XNOR2X1TH U1396 ( .A(n1110), .B(n1106), .Y(n650) );
  XNOR2X1TH U1397 ( .A(n1112), .B(n1105), .Y(n665) );
  XNOR2X1TH U1398 ( .A(n1109), .B(n1104), .Y(n685) );
  XNOR2X1TH U1399 ( .A(n1111), .B(n1104), .Y(n683) );
  XNOR2X1TH U1400 ( .A(n1115), .B(n1103), .Y(n696) );
  XNOR2X1TH U1401 ( .A(n1115), .B(n1104), .Y(n679) );
  XNOR2X1TH U1402 ( .A(n1111), .B(n1105), .Y(n666) );
  XNOR2X1TH U1403 ( .A(n1109), .B(n1105), .Y(n668) );
  XNOR2X1TH U1404 ( .A(n1111), .B(n1106), .Y(n649) );
  XNOR2X1TH U1405 ( .A(n1118), .B(n1102), .Y(n710) );
  XNOR2XLTH U1406 ( .A(n1123), .B(n1104), .Y(n687) );
  XNOR2XLTH U1407 ( .A(n1123), .B(n1105), .Y(n670) );
  XNOR2XLTH U1408 ( .A(n1123), .B(n1106), .Y(n653) );
  XNOR2XLTH U1409 ( .A(n1123), .B(n1107), .Y(n636) );
  NAND2XLTH U1410 ( .A(n1121), .B(n1100), .Y(n968) );
  XNOR2X1TH U1411 ( .A(n1113), .B(n1106), .Y(n647) );
  XNOR2X1TH U1412 ( .A(n1122), .B(n1102), .Y(n706) );
  XNOR2X1TH U1413 ( .A(n1121), .B(n1102), .Y(n707) );
  XNOR2X1TH U1414 ( .A(n1116), .B(n1104), .Y(n678) );
  XNOR2X1TH U1415 ( .A(n1118), .B(n1103), .Y(n693) );
  XNOR2X1TH U1416 ( .A(n1112), .B(n1106), .Y(n648) );
  XNOR2X1TH U1417 ( .A(n1116), .B(n1105), .Y(n661) );
  XNOR2X1TH U1418 ( .A(n1117), .B(n1104), .Y(n677) );
  XNOR2X1TH U1419 ( .A(n1110), .B(n1107), .Y(n633) );
  XNOR2X1TH U1420 ( .A(n1111), .B(n1107), .Y(n632) );
  XNOR2X1TH U1421 ( .A(n1120), .B(n1102), .Y(n708) );
  XNOR2X1TH U1422 ( .A(n1120), .B(n1103), .Y(n691) );
  XNOR2X1TH U1423 ( .A(n1122), .B(n1103), .Y(n689) );
  XNOR2X1TH U1424 ( .A(n1121), .B(n1104), .Y(n673) );
  XNOR2X1TH U1425 ( .A(n1113), .B(n1107), .Y(n630) );
  XNOR2X1TH U1426 ( .A(n1121), .B(n1103), .Y(n690) );
  XNOR2X1TH U1427 ( .A(n1118), .B(n1104), .Y(n676) );
  XNOR2X1TH U1428 ( .A(n1118), .B(n1105), .Y(n659) );
  XNOR2X1TH U1429 ( .A(n1117), .B(n1105), .Y(n660) );
  XNOR2X1TH U1430 ( .A(n1122), .B(n1104), .Y(n672) );
  XNOR2X1TH U1431 ( .A(n1118), .B(n1106), .Y(n642) );
  XNOR2X1TH U1432 ( .A(n1118), .B(n1107), .Y(n625) );
  XNOR2X1TH U1433 ( .A(n1122), .B(n1105), .Y(n655) );
  XNOR2X1TH U1434 ( .A(n1122), .B(n1106), .Y(n638) );
  XNOR2X1TH U1435 ( .A(n1122), .B(n1107), .Y(n621) );
  XOR2X1 U1436 ( .A(n341), .B(n352), .Y(n951) );
  AND2X2 U1437 ( .A(n445), .B(n929), .Y(n874) );
  OR2XLTH U1438 ( .A(n1052), .B(n1158), .Y(n889) );
  OAI22XLTH U1439 ( .A0(n712), .A1(n1051), .B0(n711), .B1(n795), .Y(n562) );
  OAI22XLTH U1440 ( .A0(n710), .A1(n795), .B0(n711), .B1(n1051), .Y(n561) );
  OAI22XLTH U1441 ( .A0(n708), .A1(n1051), .B0(n707), .B1(n795), .Y(n558) );
  OAI22XLTH U1442 ( .A0(n752), .A1(n788), .B0(n751), .B1(n1099), .Y(n603) );
  NOR2XLTH U1443 ( .A(n703), .B(n794), .Y(n1023) );
  OR2XLTH U1444 ( .A(n720), .B(n795), .Y(n882) );
  OR2XLTH U1445 ( .A(n700), .B(n794), .Y(n1045) );
  OAI22XLTH U1446 ( .A0(n706), .A1(n795), .B0(n707), .B1(n1051), .Y(n557) );
  OAI22XLTH U1447 ( .A0(n708), .A1(n795), .B0(n709), .B1(n1051), .Y(n559) );
  OAI22XLTH U1448 ( .A0(n733), .A1(n1050), .B0(n732), .B1(n796), .Y(n584) );
  OR2XLTH U1449 ( .A(n701), .B(n1053), .Y(n1044) );
  OR2XLTH U1450 ( .A(n709), .B(n795), .Y(n920) );
  OAI22XLTH U1451 ( .A0(n691), .A1(n1053), .B0(n690), .B1(n794), .Y(n540) );
  OAI22XLTH U1452 ( .A0(n691), .A1(n794), .B0(n692), .B1(n1053), .Y(n541) );
  OR2XLTH U1453 ( .A(n710), .B(n1051), .Y(n919) );
  AO21XLTH U1454 ( .A0(n1050), .A1(n796), .B0(n1160), .Y(n573) );
  AO21XLTH U1455 ( .A0(n1051), .A1(n795), .B0(n1164), .Y(n555) );
  AO21XLTH U1456 ( .A0(n1053), .A1(n794), .B0(n1163), .Y(n537) );
  AO21XLTH U1457 ( .A0(n1052), .A1(n792), .B0(n1158), .Y(n501) );
  AO21XLTH U1458 ( .A0(n1049), .A1(n791), .B0(n1157), .Y(n483) );
  AO21XLTH U1459 ( .A0(n1054), .A1(n793), .B0(n1159), .Y(n519) );
  AO21XLTH U1460 ( .A0(n788), .A1(n1099), .B0(n1165), .Y(n319) );
  ADDHX1 U1461 ( .A(n448), .B(n513), .CO(n362), .S(n363) );
  NAND2XLTH U1462 ( .A(n1153), .B(n1164), .Y(n1021) );
  OR2XLTH U1463 ( .A(n721), .B(n1051), .Y(n881) );
  OR2XLTH U1464 ( .A(n671), .B(n792), .Y(n888) );
  INVXL U1465 ( .A(n1118), .Y(n1146) );
  INVXL U1466 ( .A(n1111), .Y(n1150) );
  INVXL U1467 ( .A(n289), .Y(n1151) );
endmodule


module multiplier_0 ( data1, data2, out );
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] out;
  wire   N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, abs_data2_15_, N87, N88, N89, N90, N91, N92, N93,
         N94, N95, N96, N97, N98, N99, N100, N101, N102, n4, n12, n310, n320,
         n330, n340, n350, n360, n37, n38, n123, n124, n125, n126, n129, n2,
         n3, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17, n18, n20, n210,
         n230, n240, n250, n270, n280, n290, n300, n39, n40, n41, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n540, n550, n560, n570, n580,
         n600, n610, n620, n630, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153;
  wire   [15:0] abs_data1;
  wire   [30:15] abs_c;

  multiplier_0_DW01_inc_0 add_41 ( .A({n145, n2, n3, n146, n6, n7, n8, n9, n10, 
        n11, n13, n14, n15, n16, n17, n18}), .SUM({N102, N101, N100, N99, N98, 
        N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87}) );
  multiplier_0_DW01_inc_1 add_29 ( .A({n152, n44, n45, n46, n47, n48, n49, n50, 
        n51, n52, n53, n540, n550, n560, n570, n580}), .SUM({N69, N68, N67, 
        N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54}) );
  multiplier_0_DW01_inc_2 add_21 ( .A({n147, n20, n210, n149, n230, n240, n250, 
        n150, n270, n280, n290, n300, n39, n40, n41, n151}), .SUM({N36, N35, 
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21})
         );
  multiplier_0_DW_mult_uns_3 mult_36 ( .a({abs_data1[15:13], n129, n123, 
        abs_data1[10:7], n4, n12, abs_data1[4:0]}), .b({abs_data2_15_, n360, 
        n600, n37, n610, n330, n620, n350, n126, n340, n125, n320, n630, n310, 
        n124, n38}), .product_30_(abs_c[30]), .product_29_(abs_c[29]), 
        .product_28_(abs_c[28]), .product_27_(abs_c[27]), .product_26_(
        abs_c[26]), .product_25_(abs_c[25]), .product_24_(abs_c[24]), 
        .product_23_(abs_c[23]), .product_22_(abs_c[22]), .product_21_(
        abs_c[21]), .product_20_(abs_c[20]), .product_19_(abs_c[19]), 
        .product_18_(abs_c[18]), .product_17_(abs_c[17]), .product_16_(
        abs_c[16]), .product_15_(abs_c[15]) );
  INVX2 U2 ( .A(n135), .Y(n18) );
  BUFX8 U3 ( .A(abs_c[15]), .Y(n135) );
  OAI2B2X2TH U4 ( .A1N(N32), .A0(n147), .B0(n139), .B1(n230), .Y(n123) );
  OAI2B2X1 U5 ( .A1N(N23), .A0(n147), .B0(n139), .B1(n40), .Y(abs_data1[2]) );
  INVX6 U6 ( .A(abs_c[18]), .Y(n15) );
  INVX5 U7 ( .A(abs_c[26]), .Y(n6) );
  AO2B2X4 U8 ( .B0(N98), .B1(n142), .A0(abs_c[26]), .A1N(n141), .Y(out[11]) );
  INVX4 U9 ( .A(abs_c[24]), .Y(n8) );
  INVX4 U10 ( .A(abs_c[16]), .Y(n17) );
  INVX5 U11 ( .A(data1[11]), .Y(n230) );
  INVX6 U12 ( .A(abs_c[20]), .Y(n13) );
  INVX2 U13 ( .A(abs_c[23]), .Y(n9) );
  AO2B2X4 U14 ( .B0(N95), .B1(n142), .A0(abs_c[23]), .A1N(n140), .Y(out[8]) );
  BUFX6 U15 ( .A(abs_c[21]), .Y(n138) );
  BUFX6 U16 ( .A(abs_c[22]), .Y(n136) );
  CLKINVX2TH U17 ( .A(data1[10]), .Y(n240) );
  OAI2BB2X1TH U18 ( .B0(n14), .B1(n140), .A0N(N91), .A1N(n141), .Y(out[4]) );
  INVX1TH U19 ( .A(abs_c[25]), .Y(n7) );
  INVX18 U20 ( .A(n139), .Y(n147) );
  OAI2BB2X2TH U21 ( .B0(n146), .B1(n141), .A0N(N99), .A1N(n141), .Y(out[12])
         );
  OAI2B2XL U22 ( .A1N(N30), .A0(n147), .B0(n139), .B1(n250), .Y(abs_data1[9])
         );
  INVX4 U23 ( .A(abs_c[19]), .Y(n14) );
  INVX2 U24 ( .A(data1[0]), .Y(n151) );
  BUFX16 U25 ( .A(data1[15]), .Y(n139) );
  INVX2 U26 ( .A(abs_c[17]), .Y(n16) );
  CLKINVX1TH U27 ( .A(data1[12]), .Y(n149) );
  CLKINVX1TH U28 ( .A(data1[8]), .Y(n150) );
  OAI2BB2X2 U29 ( .B0(n145), .B1(n140), .A0N(N102), .A1N(n141), .Y(out[15]) );
  OAI2B2X1TH U30 ( .A1N(N26), .A0(n147), .B0(n139), .B1(n290), .Y(n12) );
  OAI2B2X1TH U31 ( .A1N(N22), .A0(n147), .B0(n139), .B1(n41), .Y(abs_data1[1])
         );
  INVXLTH U32 ( .A(data1[13]), .Y(n148) );
  OAI2BB2X1TH U33 ( .B0(n8), .B1(n140), .A0N(N96), .A1N(n142), .Y(out[9]) );
  OAI2BB2X2TH U34 ( .B0(n13), .B1(n140), .A0N(N92), .A1N(n141), .Y(out[5]) );
  OAI2BB2X2 U35 ( .B0(n7), .B1(n141), .A0N(N97), .A1N(n142), .Y(out[10]) );
  XNOR2XLTH U36 ( .A(n147), .B(data2[15]), .Y(n137) );
  INVX2TH U37 ( .A(abs_c[27]), .Y(n146) );
  OAI2B2X1TH U38 ( .A1N(N24), .A0(n147), .B0(n139), .B1(n39), .Y(abs_data1[3])
         );
  NOR2BXL U39 ( .AN(N36), .B(n147), .Y(abs_data1[15]) );
  INVXLTH U40 ( .A(abs_c[29]), .Y(n2) );
  INVXLTH U41 ( .A(n136), .Y(n10) );
  AO2B2XLTH U42 ( .B0(N93), .B1(n142), .A0(n138), .A1N(n140), .Y(out[6]) );
  AO2B2XLTH U43 ( .B0(N94), .B1(n142), .A0(n136), .A1N(n140), .Y(out[7]) );
  OAI2B2XL U44 ( .A1N(N21), .A0(n147), .B0(n139), .B1(n151), .Y(abs_data1[0])
         );
  OAI2B2X4 U45 ( .A1N(N31), .A0(n147), .B0(n139), .B1(n240), .Y(abs_data1[10])
         );
  CLKINVX1TH U46 ( .A(data1[9]), .Y(n250) );
  OAI2B2X4 U47 ( .A1N(N33), .A0(n147), .B0(n139), .B1(n149), .Y(n129) );
  INVX10 U48 ( .A(abs_c[28]), .Y(n3) );
  OAI2B2X4 U49 ( .A1N(N34), .A0(n147), .B0(n139), .B1(n148), .Y(abs_data1[13])
         );
  OAI2B2X2 U50 ( .A1N(N35), .A0(n147), .B0(n139), .B1(n20), .Y(abs_data1[14])
         );
  INVXLTH U51 ( .A(data1[3]), .Y(n39) );
  INVXLTH U52 ( .A(data1[2]), .Y(n40) );
  INVXLTH U53 ( .A(data1[6]), .Y(n280) );
  INVXLTH U54 ( .A(data1[4]), .Y(n300) );
  INVXLTH U55 ( .A(data1[1]), .Y(n41) );
  INVXLTH U56 ( .A(data1[5]), .Y(n290) );
  INVXLTH U57 ( .A(data2[4]), .Y(n540) );
  INVXLTH U58 ( .A(data2[8]), .Y(n50) );
  INVXLTH U59 ( .A(data1[7]), .Y(n270) );
  INVXLTH U60 ( .A(data2[5]), .Y(n53) );
  INVXLTH U61 ( .A(data2[7]), .Y(n51) );
  INVXLTH U62 ( .A(data2[6]), .Y(n52) );
  INVXLTH U63 ( .A(data2[12]), .Y(n46) );
  INVXLTH U64 ( .A(data2[9]), .Y(n49) );
  INVXLTH U65 ( .A(data2[10]), .Y(n48) );
  INVXLTH U66 ( .A(data2[11]), .Y(n47) );
  INVXLTH U67 ( .A(data2[3]), .Y(n550) );
  INVXLTH U68 ( .A(data2[2]), .Y(n560) );
  INVXLTH U69 ( .A(data2[14]), .Y(n44) );
  INVXLTH U70 ( .A(data2[13]), .Y(n45) );
  CLKINVX1TH U71 ( .A(data1[14]), .Y(n20) );
  INVXLTH U72 ( .A(data1[13]), .Y(n210) );
  INVXLTH U73 ( .A(data2[0]), .Y(n580) );
  INVXLTH U74 ( .A(data2[1]), .Y(n570) );
  INVX4TH U75 ( .A(data2[15]), .Y(n152) );
  OAI2B2X1TH U76 ( .A1N(N68), .A0(n152), .B0(data2[15]), .B1(n44), .Y(n360) );
  OAI2B2X1TH U77 ( .A1N(N58), .A0(n152), .B0(data2[15]), .B1(n540), .Y(n320)
         );
  OAI2B2X1TH U78 ( .A1N(N62), .A0(n152), .B0(data2[15]), .B1(n50), .Y(n350) );
  OAI2B2XLTH U79 ( .A1N(N59), .A0(n152), .B0(data2[15]), .B1(n53), .Y(n125) );
  OAI2B2XLTH U80 ( .A1N(N61), .A0(n152), .B0(data2[15]), .B1(n51), .Y(n126) );
  OAI2B2X1TH U81 ( .A1N(N60), .A0(n152), .B0(data2[15]), .B1(n52), .Y(n340) );
  OAI2B2X1TH U82 ( .A1N(N66), .A0(n152), .B0(data2[15]), .B1(n46), .Y(n37) );
  OAI2B2XLTH U83 ( .A1N(N63), .A0(n152), .B0(data2[15]), .B1(n49), .Y(n620) );
  OAI2B2X1TH U84 ( .A1N(N64), .A0(n152), .B0(data2[15]), .B1(n48), .Y(n330) );
  OAI2B2XLTH U85 ( .A1N(N65), .A0(n152), .B0(data2[15]), .B1(n47), .Y(n610) );
  OAI2B2XLTH U86 ( .A1N(N57), .A0(n152), .B0(data2[15]), .B1(n550), .Y(n630)
         );
  OAI2B2X1TH U87 ( .A1N(N56), .A0(n152), .B0(data2[15]), .B1(n560), .Y(n310)
         );
  NOR2BXLTH U88 ( .AN(N69), .B(n152), .Y(abs_data2_15_) );
  OAI2B2XLTH U89 ( .A1N(N67), .A0(n152), .B0(data2[15]), .B1(n45), .Y(n600) );
  OAI2B2X1TH U90 ( .A1N(N54), .A0(n152), .B0(data2[15]), .B1(n153), .Y(n38) );
  INVXLTH U91 ( .A(data2[0]), .Y(n153) );
  OAI2B2XLTH U92 ( .A1N(N55), .A0(n152), .B0(data2[15]), .B1(n570), .Y(n124)
         );
  INVXLTH U93 ( .A(n138), .Y(n11) );
  INVXLTH U94 ( .A(abs_c[30]), .Y(n145) );
  CLKBUFX1TH U95 ( .A(n137), .Y(n143) );
  BUFX3TH U96 ( .A(n143), .Y(n140) );
  CLKBUFX2TH U97 ( .A(n143), .Y(n142) );
  BUFX3TH U98 ( .A(n143), .Y(n141) );
  OAI2BB2XLTH U99 ( .B0(n144), .B1(n141), .A0N(N87), .A1N(n142), .Y(out[0]) );
  AO2B2X4 U100 ( .B0(N101), .B1(n141), .A0(abs_c[29]), .A1N(n140), .Y(out[14])
         );
  OAI2B2XLTH U101 ( .A1N(N27), .A0(n147), .B0(n139), .B1(n280), .Y(n4) );
  OAI2B2X1 U102 ( .A1N(N25), .A0(n147), .B0(n139), .B1(n300), .Y(abs_data1[4])
         );
  OAI2B2XLTH U103 ( .A1N(N28), .A0(n147), .B0(n139), .B1(n270), .Y(
        abs_data1[7]) );
  OAI2B2XLTH U104 ( .A1N(N29), .A0(n147), .B0(n139), .B1(n150), .Y(
        abs_data1[8]) );
  AO2B2X4 U105 ( .B0(N100), .B1(n141), .A0(abs_c[28]), .A1N(n140), .Y(out[13])
         );
  OAI2BB2XLTH U106 ( .B0(n17), .B1(n140), .A0N(N88), .A1N(n141), .Y(out[1]) );
  OAI2BB2XLTH U107 ( .B0(n16), .B1(n140), .A0N(N89), .A1N(n141), .Y(out[2]) );
  OAI2BB2XLTH U108 ( .B0(n15), .B1(n140), .A0N(N90), .A1N(n141), .Y(out[3]) );
  INVXLTH U109 ( .A(n135), .Y(n144) );
endmodule


module bpsk_adder ( out_b, in1, in2 );
  output [15:0] out_b;
  input [11:0] in1;
  input in2;
  wire   n62, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n39, n40, n43, n44,
         n45, n46, n47, n48, n61;

  OAI21BX4 U3 ( .A0(n39), .A1(n5), .B0N(n6), .Y(n62) );
  BUFX2 U4 ( .A(in1[6]), .Y(out_b[6]) );
  NAND2X2 U5 ( .A(in1[10]), .B(n45), .Y(n46) );
  INVX4 U6 ( .A(n13), .Y(n45) );
  BUFX6 U7 ( .A(n4), .Y(n39) );
  NOR2XL U8 ( .A(n40), .B(n44), .Y(n4) );
  CLKNAND2X8 U9 ( .A(n46), .B(n47), .Y(out_b[10]) );
  XOR2X3 U10 ( .A(in2), .B(in1[9]), .Y(n13) );
  CLKBUFX16 U11 ( .A(in1[2]), .Y(out_b[2]) );
  CLKBUFX16 U12 ( .A(in1[5]), .Y(out_b[5]) );
  NAND2X2TH U13 ( .A(n43), .B(n8), .Y(out_b[11]) );
  BUFX10 U14 ( .A(n62), .Y(out_b[12]) );
  BUFX2TH U15 ( .A(out_b[12]), .Y(out_b[14]) );
  CLKBUFX2TH U16 ( .A(in1[8]), .Y(out_b[8]) );
  OR2XLTH U17 ( .A(in2), .B(out_b[9]), .Y(n40) );
  CLKBUFX16 U18 ( .A(in1[0]), .Y(out_b[0]) );
  INVX4TH U19 ( .A(in1[9]), .Y(out_b[9]) );
  CLKNAND2X4 U20 ( .A(n44), .B(n13), .Y(n47) );
  OR3X2 U21 ( .A(in1[7]), .B(in1[0]), .C(out_b[8]), .Y(n12) );
  CLKBUFX1TH U22 ( .A(in1[1]), .Y(out_b[1]) );
  AOI222XL U23 ( .A0(in2), .A1(in1[9]), .B0(n44), .B1(n61), .C0(in1[10]), .C1(
        out_b[9]), .Y(n7) );
  INVX2TH U24 ( .A(in1[10]), .Y(n44) );
  CLKNAND2X8 U25 ( .A(n48), .B(in1[11]), .Y(n5) );
  BUFX2TH U26 ( .A(out_b[12]), .Y(out_b[13]) );
  OAI21X1 U27 ( .A0(n39), .A1(n6), .B0(n5), .Y(n8) );
  BUFX3TH U28 ( .A(in1[4]), .Y(out_b[4]) );
  BUFX3TH U29 ( .A(in1[3]), .Y(out_b[3]) );
  INVXLTH U30 ( .A(in2), .Y(n61) );
  OR2XL U31 ( .A(n7), .B(n5), .Y(n43) );
  OR3X2 U32 ( .A(n9), .B(n10), .C(n11), .Y(n48) );
  BUFX20 U33 ( .A(in1[7]), .Y(out_b[7]) );
  OR3XLTH U34 ( .A(n12), .B(in1[5]), .C(in1[6]), .Y(n9) );
  OR3XLTH U35 ( .A(in1[2]), .B(in1[3]), .C(in1[1]), .Y(n11) );
  BUFX2TH U36 ( .A(out_b[12]), .Y(out_b[15]) );
  NOR3X1TH U37 ( .A(in1[10]), .B(in1[9]), .C(n61), .Y(n6) );
  OR3XLTH U38 ( .A(in1[10]), .B(in1[9]), .C(in1[4]), .Y(n10) );
endmodule


module qu_table_tc_test_1 ( out, in, clk, reset, test_si, test_se );
  output [4:0] out;
  input [15:0] in;
  input clk, reset, test_si, test_se;
  wire   n321, n322, n324, n325, n225, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n300, n301;

  NOR4X2 U33 ( .A(n288), .B(in[7]), .C(n71), .D(n73), .Y(n93) );
  OAI31X1 U109 ( .A0(n102), .A1(in[7]), .A2(n103), .B0(n74), .Y(n101) );
  NOR3X1 U110 ( .A(n294), .B(n297), .C(n296), .Y(n103) );
  OAI31X1 U122 ( .A0(in[11]), .A1(in[13]), .A2(in[12]), .B0(n110), .Y(n116) );
  NOR3X1 U133 ( .A(n240), .B(n244), .C(n279), .Y(n133) );
  SDFFRQXLTH out_reg_1_ ( .D(n322), .SI(out[0]), .SE(n301), .CK(clk), .RN(n257), .Q(out[1]) );
  SDFFRQXLTH out_reg_4_ ( .D(n325), .SI(out[3]), .SE(n300), .CK(clk), .RN(n257), .Q(out[4]) );
  SDFFRQXLTH out_reg_3_ ( .D(n324), .SI(out[2]), .SE(n300), .CK(clk), .RN(
        reset), .Q(out[3]) );
  SDFFRQXLTH out_reg_0_ ( .D(n321), .SI(test_si), .SE(n301), .CK(clk), .RN(
        n257), .Q(out[0]) );
  SDFFRQXLTH out_reg_2_ ( .D(n225), .SI(out[1]), .SE(n301), .CK(clk), .RN(n257), .Q(out[2]) );
  AOI2BB1X1 U3 ( .A0N(n92), .A1N(n291), .B0(n288), .Y(n71) );
  INVX2 U4 ( .A(n110), .Y(n288) );
  AOI21X1TH U5 ( .A0(n55), .A1(n122), .B0(n137), .Y(n136) );
  BUFX10 U6 ( .A(n113), .Y(n236) );
  NOR4X1 U7 ( .A(n56), .B(n57), .C(n36), .D(n282), .Y(n43) );
  BUFX20 U8 ( .A(n120), .Y(n237) );
  BUFX10 U9 ( .A(n50), .Y(n238) );
  OAI21X1 U10 ( .A0(n90), .A1(n253), .B0(n91), .Y(n62) );
  NOR4X6 U11 ( .A(in[11]), .B(in[12]), .C(in[13]), .D(in[14]), .Y(n91) );
  NOR3X6 U12 ( .A(n236), .B(n249), .C(n46), .Y(n75) );
  INVX4 U13 ( .A(n91), .Y(n284) );
  CLKXOR2X2 U14 ( .A(n144), .B(n291), .Y(n53) );
  NAND2X1 U15 ( .A(n145), .B(n292), .Y(n144) );
  BUFX4 U16 ( .A(n119), .Y(n239) );
  NOR2BX8 U17 ( .AN(n238), .B(n38), .Y(n121) );
  AOI31X1 U18 ( .A0(n251), .A1(n275), .A2(n81), .B0(n270), .Y(n77) );
  INVX1 U19 ( .A(n130), .Y(n275) );
  NOR2BX8 U20 ( .AN(n122), .B(n251), .Y(n86) );
  NAND3X4 U21 ( .A(n138), .B(n273), .C(n139), .Y(n122) );
  OAI32X2 U22 ( .A0(n36), .A1(in[15]), .A2(n281), .B0(n37), .B1(n286), .Y(n324) );
  NAND2X8 U23 ( .A(n108), .B(n104), .Y(n126) );
  XOR2X8 U24 ( .A(n108), .B(n296), .Y(n127) );
  NAND2X4 U25 ( .A(n297), .B(n280), .Y(n108) );
  OAI31X4 U26 ( .A0(n82), .A1(n237), .A2(n53), .B0(n134), .Y(n113) );
  AOI31X1 U27 ( .A0(n272), .A1(n55), .A2(n135), .B0(n269), .Y(n134) );
  BUFX8 U28 ( .A(n40), .Y(n249) );
  INVXLTH U29 ( .A(in[1]), .Y(n297) );
  NAND2X4 U30 ( .A(n255), .B(n256), .Y(n115) );
  CLKNAND2X2 U31 ( .A(in[10]), .B(n254), .Y(n255) );
  CLKINVX2TH U32 ( .A(in[6]), .Y(n293) );
  CLKBUFX2TH U34 ( .A(n80), .Y(n251) );
  NAND3XL U35 ( .A(n55), .B(n53), .C(n86), .Y(n54) );
  CLKINVX1TH U36 ( .A(n62), .Y(n271) );
  AOI32X2 U37 ( .A0(n245), .A1(n59), .A2(n65), .B0(n66), .B1(n286), .Y(n63) );
  NAND4X2 U38 ( .A(n67), .B(n68), .C(n58), .D(n69), .Y(n66) );
  NOR4BX4 U39 ( .AN(n67), .B(n88), .C(n89), .D(n62), .Y(n87) );
  NOR2X8 U40 ( .A(n108), .B(in[2]), .Y(n150) );
  NOR2X8 U41 ( .A(n149), .B(in[4]), .Y(n148) );
  NAND2X6 U42 ( .A(n150), .B(n295), .Y(n149) );
  NOR2X8 U43 ( .A(n146), .B(in[6]), .Y(n145) );
  NAND2X8 U44 ( .A(n148), .B(n294), .Y(n146) );
  NAND2X4 U45 ( .A(n253), .B(n142), .Y(n256) );
  INVX2 U46 ( .A(n142), .Y(n254) );
  INVX10 U47 ( .A(n53), .Y(n277) );
  NOR2XL U48 ( .A(n292), .B(n293), .Y(n70) );
  BUFX10 U49 ( .A(n123), .Y(n242) );
  NAND2X2 U50 ( .A(n293), .B(n105), .Y(n102) );
  NOR2X2 U51 ( .A(in[9]), .B(n143), .Y(n142) );
  BUFX3 U52 ( .A(n126), .Y(n244) );
  AOI21X1TH U53 ( .A0(n294), .A1(n106), .B0(n293), .Y(n73) );
  OAI21BX1TH U54 ( .A0(n129), .A1(n131), .B0N(n239), .Y(n47) );
  AOI21XLTH U55 ( .A0(n242), .A1(n278), .B0(n130), .Y(n137) );
  CLKBUFX3 U56 ( .A(n94), .Y(n243) );
  NAND3X2TH U57 ( .A(n294), .B(n293), .C(n107), .Y(n72) );
  OAI21X2 U58 ( .A0(n70), .A1(n287), .B0(n71), .Y(n58) );
  NAND2X2 U59 ( .A(n241), .B(n101), .Y(n61) );
  INVX2 U60 ( .A(n69), .Y(n282) );
  AND4X1TH U61 ( .A(n109), .B(n289), .C(n42), .D(n253), .Y(n36) );
  NAND3XL U62 ( .A(n53), .B(n54), .C(n55), .Y(n34) );
  OAI221XL U63 ( .A0(n59), .A1(n287), .B0(n60), .B1(n61), .C0(n271), .Y(n56)
         );
  BUFX8 U64 ( .A(n127), .Y(n240) );
  OAI31X2 U65 ( .A0(n85), .A1(n133), .A2(n251), .B0(n277), .Y(n132) );
  INVX18 U66 ( .A(n251), .Y(n278) );
  NOR4BX4 U67 ( .AN(n82), .B(n275), .C(n277), .D(n251), .Y(n114) );
  CLKNAND2X2 U68 ( .A(in[1]), .B(in[0]), .Y(n104) );
  NOR2X2 U69 ( .A(n284), .B(in[10]), .Y(n99) );
  NOR4X1 U70 ( .A(n38), .B(n39), .C(n249), .D(n41), .Y(n37) );
  OAI211X4 U71 ( .A0(n114), .A1(n115), .B0(n116), .C0(n117), .Y(n46) );
  AOI22XL U72 ( .A0(n118), .A1(n288), .B0(in[14]), .B1(n285), .Y(n117) );
  CLKXOR2X4 U73 ( .A(n143), .B(n290), .Y(n130) );
  CLKINVX12 U74 ( .A(in[8]), .Y(n291) );
  NOR2X2TH U75 ( .A(n294), .B(n246), .Y(n247) );
  AND4X2TH U76 ( .A(n75), .B(n76), .C(n77), .D(n52), .Y(n35) );
  NAND3X2 U77 ( .A(n237), .B(n274), .C(n136), .Y(n51) );
  INVXLTH U78 ( .A(n51), .Y(n269) );
  INVX2TH U79 ( .A(in[9]), .Y(n290) );
  XOR2XLTH U80 ( .A(n145), .B(n292), .Y(n80) );
  NAND2X2TH U81 ( .A(n242), .B(n141), .Y(n85) );
  INVXLTH U82 ( .A(n74), .Y(n289) );
  AOI31X1TH U83 ( .A0(n75), .A1(n268), .A2(in[15]), .B0(n87), .Y(n225) );
  OAI21X3TH U84 ( .A0(n35), .A1(n286), .B0(n63), .Y(n321) );
  NOR3BX1TH U85 ( .AN(n34), .B(n45), .C(n41), .Y(n44) );
  NOR2X1TH U86 ( .A(n288), .B(in[8]), .Y(n65) );
  NAND3X1 U87 ( .A(in[12]), .B(in[11]), .C(in[14]), .Y(n118) );
  BUFX5 U88 ( .A(n99), .Y(n241) );
  NOR4BX4 U89 ( .AN(n72), .B(n98), .C(n284), .D(n73), .Y(n97) );
  XOR2XL U90 ( .A(n146), .B(n293), .Y(n123) );
  NAND3X4 U91 ( .A(n59), .B(n61), .C(n241), .Y(n69) );
  CLKINVX4 U92 ( .A(in[10]), .Y(n253) );
  NAND2BX8 U93 ( .AN(n144), .B(n291), .Y(n143) );
  NAND4BX2 U94 ( .AN(n46), .B(n47), .C(n48), .D(n49), .Y(n41) );
  NOR3X6 U95 ( .A(n36), .B(n95), .C(n96), .Y(n67) );
  XOR2X8 U96 ( .A(n148), .B(n294), .Y(n138) );
  INVX6 U97 ( .A(in[5]), .Y(n294) );
  NOR2X5TH U98 ( .A(n252), .B(n55), .Y(n129) );
  NOR3X2 U99 ( .A(n82), .B(n130), .C(n278), .Y(n131) );
  CLKINVX1TH U100 ( .A(in[3]), .Y(n295) );
  INVXLTH U101 ( .A(in[0]), .Y(n280) );
  CLKINVX1TH U102 ( .A(n138), .Y(n279) );
  INVXLTH U103 ( .A(n242), .Y(n273) );
  INVX3TH U104 ( .A(n115), .Y(n276) );
  NAND3XLTH U105 ( .A(n291), .B(n290), .C(n292), .Y(n98) );
  INVXLTH U106 ( .A(n49), .Y(n270) );
  AOI31X4TH U107 ( .A0(n33), .A1(n34), .A2(n35), .B0(n286), .Y(n325) );
  CLKINVX1TH U108 ( .A(n258), .Y(n257) );
  NAND3XLTH U111 ( .A(n238), .B(n51), .C(n52), .Y(n45) );
  NOR2X2TH U112 ( .A(in[10]), .B(in[9]), .Y(n110) );
  OAI21XLTH U113 ( .A0(in[6]), .A1(in[7]), .B0(in[9]), .Y(n109) );
  OR2XLTH U114 ( .A(n247), .B(n102), .Y(n245) );
  OR2XLTH U115 ( .A(n104), .B(n296), .Y(n246) );
  CLKINVX1TH U116 ( .A(in[2]), .Y(n296) );
  NOR2BX2TH U117 ( .AN(n100), .B(in[7]), .Y(n59) );
  NOR3X4TH U118 ( .A(n78), .B(n86), .C(n274), .Y(n38) );
  OAI21XLTH U119 ( .A0(n78), .A1(n277), .B0(n79), .Y(n52) );
  NOR2X1TH U120 ( .A(n278), .B(n242), .Y(n78) );
  NAND3X3 U123 ( .A(n115), .B(n239), .C(n86), .Y(n49) );
  OAI21X6 U124 ( .A0(n278), .A1(n53), .B0(n55), .Y(n120) );
  NOR3BX4 U125 ( .AN(n47), .B(n39), .C(n112), .Y(n33) );
  OAI21XL U126 ( .A0(n130), .A1(n132), .B0(n115), .Y(n119) );
  AND3X2 U127 ( .A(n92), .B(n290), .C(n291), .Y(n90) );
  NOR2X8 U128 ( .A(n290), .B(n291), .Y(n74) );
  AOI21X4 U129 ( .A0(n83), .A1(n277), .B0(n237), .Y(n79) );
  AOI211X2 U130 ( .A0(n278), .A1(n242), .B0(n129), .C0(n130), .Y(n39) );
  AND2XL U131 ( .A(n115), .B(n53), .Y(n252) );
  OAI22X2 U132 ( .A0(in[15]), .A1(n43), .B0(n44), .B1(n286), .Y(n322) );
  INVX2TH U134 ( .A(n245), .Y(n283) );
  NOR4X1 U135 ( .A(n71), .B(n93), .C(n89), .D(n288), .Y(n95) );
  INVX2TH U136 ( .A(n65), .Y(n287) );
  INVXLTH U137 ( .A(in[13]), .Y(n285) );
  NOR3X4TH U138 ( .A(n279), .B(n240), .C(n140), .Y(n84) );
  OAI21X2TH U139 ( .A0(n147), .A1(n138), .B0(n273), .Y(n82) );
  AOI211XLTH U140 ( .A0(n244), .A1(n280), .B0(n240), .C0(n128), .Y(n124) );
  NAND3X1TH U141 ( .A(in[4]), .B(in[6]), .C(n111), .Y(n100) );
  INVXLTH U142 ( .A(n112), .Y(n268) );
  INVXLTH U143 ( .A(reset), .Y(n258) );
  INVXLTH U144 ( .A(n42), .Y(n281) );
  CLKXOR2X2 U145 ( .A(n150), .B(in[3]), .Y(n128) );
  OAI31X2 U146 ( .A0(n100), .A1(n291), .A2(n292), .B0(n110), .Y(n42) );
  XNOR2X2 U147 ( .A(n149), .B(in[4]), .Y(n125) );
  OA21X2 U148 ( .A0(n84), .A1(n85), .B0(n237), .Y(n250) );
  NAND2X1TH U149 ( .A(n250), .B(n55), .Y(n50) );
  NOR2X8 U150 ( .A(n275), .B(n276), .Y(n55) );
  INVX6 U151 ( .A(n129), .Y(n274) );
  NOR3X1 U152 ( .A(n291), .B(n283), .C(n292), .Y(n89) );
  CLKINVX32 U153 ( .A(in[7]), .Y(n292) );
  NOR2XLTH U154 ( .A(n72), .B(in[7]), .Y(n92) );
  NAND2BXLTH U155 ( .AN(n244), .B(in[0]), .Y(n140) );
  AOI211XLTH U156 ( .A0(n240), .A1(n244), .B0(n128), .C0(n125), .Y(n147) );
  AOI21XLTH U157 ( .A0(in[7]), .A1(n73), .B0(n74), .Y(n60) );
  OAI211X4 U158 ( .A0(n79), .A1(n237), .B0(n48), .C0(n121), .Y(n112) );
  NOR2BXLTH U159 ( .AN(n237), .B(n84), .Y(n135) );
  NOR4BX4 U160 ( .AN(n33), .B(n236), .C(n79), .D(n270), .Y(n40) );
  AOI31XLTH U161 ( .A0(in[2]), .A1(n108), .A2(in[3]), .B0(in[4]), .Y(n107) );
  OAI21XLTH U162 ( .A0(in[3]), .A1(in[4]), .B0(in[5]), .Y(n105) );
  OAI211XLTH U163 ( .A0(in[1]), .A1(in[2]), .B0(in[4]), .C0(in[3]), .Y(n106)
         );
  NAND4XLTH U164 ( .A(n60), .B(in[7]), .C(in[9]), .D(n72), .Y(n68) );
  NOR4BX4 U165 ( .AN(n61), .B(n282), .C(n243), .D(n97), .Y(n96) );
  OR3XLTH U166 ( .A(n93), .B(in[15]), .C(n243), .Y(n88) );
  NAND2XLTH U167 ( .A(n276), .B(n83), .Y(n48) );
  OAI31XLTH U168 ( .A0(n42), .A1(n283), .A2(n292), .B0(n58), .Y(n57) );
  INVX2 U169 ( .A(in[15]), .Y(n286) );
  NOR4BX4 U170 ( .AN(n241), .B(n289), .C(n70), .D(n59), .Y(n94) );
  AOI31XLTH U171 ( .A0(n240), .A1(n140), .A2(n128), .B0(n125), .Y(n139) );
  OAI2BB1XLTH U172 ( .A0N(n128), .A1N(n125), .B0(n138), .Y(n141) );
  NAND4BX2TH U173 ( .AN(n124), .B(n125), .C(n242), .D(n279), .Y(n83) );
  AOI31XLTH U174 ( .A0(n296), .A1(n295), .A2(n104), .B0(n294), .Y(n111) );
  OAI21BXLTH U175 ( .A0(n84), .A1(n85), .B0N(n54), .Y(n76) );
  AND3XLTH U176 ( .A(n82), .B(n274), .C(n83), .Y(n81) );
  INVXL U186 ( .A(n85), .Y(n272) );
  DLY1X1TH U187 ( .A(n301), .Y(n300) );
  DLY1X1TH U188 ( .A(test_se), .Y(n301) );
endmodule


module uniform_10_test_1 ( clk, reset, out, test_si, test_se );
  output [9:0] out;
  input clk, reset, test_si, test_se;
  wire   N0, N1, N2, n3, n4, n27, n28, n29, n30, n31, n32, n33, n34;

  SDFFRQX1TH register_reg_7_ ( .D(N0), .SI(out[6]), .SE(n33), .CK(clk), .RN(n3), .Q(out[7]) );
  SDFFRQX1TH register_reg_1_ ( .D(N2), .SI(out[0]), .SE(n31), .CK(clk), .RN(n3), .Q(out[1]) );
  SDFFRQX1TH register_reg_2_ ( .D(N1), .SI(out[1]), .SE(n32), .CK(clk), .RN(n3), .Q(out[2]) );
  SDFFRQX1TH register_reg_9_ ( .D(out[0]), .SI(out[8]), .SE(n28), .CK(clk), 
        .RN(n3), .Q(out[9]) );
  SDFFRQX1TH register_reg_6_ ( .D(out[7]), .SI(out[5]), .SE(n31), .CK(clk), 
        .RN(n3), .Q(out[6]) );
  SDFFRQX1TH register_reg_5_ ( .D(out[6]), .SI(out[4]), .SE(n32), .CK(clk), 
        .RN(n3), .Q(out[5]) );
  SDFFRQX1TH register_reg_4_ ( .D(out[5]), .SI(out[3]), .SE(n34), .CK(clk), 
        .RN(n3), .Q(out[4]) );
  SDFFRQX1TH register_reg_8_ ( .D(out[9]), .SI(out[7]), .SE(n34), .CK(clk), 
        .RN(n3), .Q(out[8]) );
  SDFFRQX1TH register_reg_3_ ( .D(out[4]), .SI(out[2]), .SE(n33), .CK(clk), 
        .RN(n3), .Q(out[3]) );
  SDFFSQX2TH register_reg_0_ ( .D(out[1]), .SI(test_si), .SE(n28), .CK(clk), 
        .SN(n3), .Q(out[0]) );
  XOR2XLTH U3 ( .A(out[3]), .B(out[0]), .Y(N1) );
  XOR2XLTH U4 ( .A(out[2]), .B(out[0]), .Y(N2) );
  CLKINVX3TH U5 ( .A(n4), .Y(n3) );
  INVXLTH U6 ( .A(reset), .Y(n4) );
  XOR2XLTH U7 ( .A(out[8]), .B(out[0]), .Y(N0) );
  DLY1X1TH U28 ( .A(n29), .Y(n27) );
  INVXLTH U29 ( .A(n27), .Y(n28) );
  INVXLTH U30 ( .A(test_se), .Y(n29) );
  INVXLTH U31 ( .A(test_se), .Y(n30) );
  INVXLTH U32 ( .A(n27), .Y(n31) );
  INVXLTH U33 ( .A(n27), .Y(n32) );
  INVXLTH U34 ( .A(n30), .Y(n33) );
  INVXLTH U35 ( .A(n30), .Y(n34) );
endmodule


module uniform_10b_test_1 ( clk, reset, out, test_si, test_se );
  output [9:0] out;
  input clk, reset, test_si, test_se;
  wire   N0, N1, N2, N3, N4, N5, N6, n28, n60, n7, n31, n32, n33, n34, n35,
         n36, n37, n38;

  SDFFSQXLTH register_reg_0_ ( .D(out[1]), .SI(test_si), .SE(n32), .CK(clk), 
        .SN(n60), .Q(n28) );
  SDFFRQX1TH register_reg_2_ ( .D(N6), .SI(out[1]), .SE(n35), .CK(clk), .RN(
        n60), .Q(out[2]) );
  SDFFRQX1TH register_reg_9_ ( .D(out[0]), .SI(out[8]), .SE(n32), .CK(clk), 
        .RN(n60), .Q(out[9]) );
  SDFFRQX1TH register_reg_8_ ( .D(N0), .SI(out[7]), .SE(n38), .CK(clk), .RN(
        n60), .Q(out[8]) );
  SDFFRQX1TH register_reg_7_ ( .D(N1), .SI(out[6]), .SE(n37), .CK(clk), .RN(
        n60), .Q(out[7]) );
  SDFFRQX1TH register_reg_6_ ( .D(N2), .SI(out[5]), .SE(n36), .CK(clk), .RN(
        n60), .Q(out[6]) );
  SDFFRQX1TH register_reg_5_ ( .D(N3), .SI(out[4]), .SE(n36), .CK(clk), .RN(
        n60), .Q(out[5]) );
  SDFFRQX1TH register_reg_4_ ( .D(N4), .SI(out[3]), .SE(n38), .CK(clk), .RN(
        n60), .Q(out[4]) );
  SDFFRQX1TH register_reg_3_ ( .D(N5), .SI(out[2]), .SE(n37), .CK(clk), .RN(
        n60), .Q(out[3]) );
  SDFFRQX1TH register_reg_1_ ( .D(out[2]), .SI(out[0]), .SE(n35), .CK(clk), 
        .RN(n60), .Q(out[1]) );
  CLKINVX3TH U3 ( .A(n7), .Y(n60) );
  INVXLTH U4 ( .A(reset), .Y(n7) );
  CLKBUFX3TH U5 ( .A(n28), .Y(out[0]) );
  XOR2XLTH U6 ( .A(out[3]), .B(out[0]), .Y(N6) );
  XOR2XLTH U7 ( .A(out[4]), .B(out[0]), .Y(N5) );
  XOR2XLTH U8 ( .A(out[5]), .B(out[0]), .Y(N4) );
  XOR2XLTH U9 ( .A(out[6]), .B(out[0]), .Y(N3) );
  XOR2XLTH U10 ( .A(out[7]), .B(out[0]), .Y(N2) );
  XOR2XLTH U11 ( .A(out[8]), .B(out[0]), .Y(N1) );
  XOR2XLTH U12 ( .A(out[9]), .B(out[0]), .Y(N0) );
  DLY1X1TH U33 ( .A(n33), .Y(n31) );
  INVXLTH U34 ( .A(n31), .Y(n32) );
  INVXLTH U35 ( .A(test_se), .Y(n33) );
  INVXLTH U36 ( .A(test_se), .Y(n34) );
  INVXLTH U37 ( .A(n31), .Y(n35) );
  INVXLTH U38 ( .A(n31), .Y(n36) );
  INVXLTH U39 ( .A(n34), .Y(n37) );
  INVXLTH U40 ( .A(n34), .Y(n38) );
endmodule


module awgn_test_1 ( clk, reset, db, qu_llr, codeword, test_si, test_so, 
        test_se );
  input [2:0] db;
  output [4:0] qu_llr;
  input clk, reset, codeword, test_si, test_se;
  output test_so;
  wire   tmp2_8_, tmp2_7_, tmp2_6_, tmp2_5_, tmp2_4_, tmp2_3_, tmp2_2_,
         tmp2_1_, tmp2_0_, n3, n4, n5, n8, n9, n10;
  wire   [9:0] tmp1;
  wire   [15:0] data1;
  wire   [15:0] data2;
  wire   [15:0] segma;
  wire   [15:0] tmp;
  wire   [15:4] tmp3;
  wire   [15:0] out_n;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5;

  nco_table_log log ( .Q(data1), .A(tmp1), .CLK(clk), .CEN(1'b0) );
  nco_table_cos cos ( .Q(data2), .A({test_so, tmp2_8_, tmp2_7_, tmp2_6_, 
        tmp2_5_, tmp2_4_, tmp2_3_, tmp2_2_, tmp2_1_, tmp2_0_}), .CLK(clk), 
        .CEN(1'b0) );
  uniform_10_test_1 u ( .clk(clk), .reset(n4), .out(tmp1), .test_si(qu_llr[4]), 
        .test_se(n9) );
  uniform_10b_test_1 v ( .clk(clk), .reset(n4), .out({test_so, tmp2_8_, 
        tmp2_7_, tmp2_6_, tmp2_5_, tmp2_4_, tmp2_3_, tmp2_2_, tmp2_1_, tmp2_0_}), .test_si(tmp1[9]), .test_se(n10) );
  segma_table s1 ( .out({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        segma[13:0]}), .in(db) );
  multiplier_1 m0 ( .data1(data1), .data2(data2), .out(tmp) );
  multiplier_0 m1 ( .data1(tmp), .data2({1'b0, 1'b1, segma[13:0]}), .out({tmp3, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5}) );
  bpsk_adder b0 ( .out_b(out_n), .in1(tmp3), .in2(codeword) );
  qu_table_tc_test_1 q2 ( .out(qu_llr), .in({out_n[15:14], n3, out_n[12:0]}), 
        .clk(clk), .reset(n4), .test_si(test_si), .test_se(test_se) );
  BUFX4 U2 ( .A(out_n[13]), .Y(n3) );
  CLKINVX1TH U3 ( .A(n5), .Y(n4) );
  INVXLTH U6 ( .A(reset), .Y(n5) );
  INVXLTH U7 ( .A(test_se), .Y(n8) );
  INVXLTH U8 ( .A(n8), .Y(n9) );
  INVXLTH U9 ( .A(n8), .Y(n10) );
endmodule


module SIPO_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  ADDHXLTH U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXLTH U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXLTH U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXLTH U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXLTH U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXLTH U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXLTH U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXLTH U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVXLTH U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2XLTH U2 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
endmodule


module SIPO_DW01_inc_1 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  ADDHXLTH U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXLTH U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXLTH U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXLTH U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXLTH U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXLTH U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXLTH U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXLTH U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  INVXLTH U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2XLTH U2 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
endmodule


module SIPO_test_1 ( out0, out1, out2, out3, out4, out5, out6, out7, out8, 
        out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, 
        out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, 
        out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, 
        out39, out40, out41, out42, out43, out44, out45, out46, out47, count1, 
        count2, in, reset, clk, test_si, test_se );
  output [4:0] out0;
  output [4:0] out1;
  output [4:0] out2;
  output [4:0] out3;
  output [4:0] out4;
  output [4:0] out5;
  output [4:0] out6;
  output [4:0] out7;
  output [4:0] out8;
  output [4:0] out9;
  output [4:0] out10;
  output [4:0] out11;
  output [4:0] out12;
  output [4:0] out13;
  output [4:0] out14;
  output [4:0] out15;
  output [4:0] out16;
  output [4:0] out17;
  output [4:0] out18;
  output [4:0] out19;
  output [4:0] out20;
  output [4:0] out21;
  output [4:0] out22;
  output [4:0] out23;
  output [4:0] out24;
  output [4:0] out25;
  output [4:0] out26;
  output [4:0] out27;
  output [4:0] out28;
  output [4:0] out29;
  output [4:0] out30;
  output [4:0] out31;
  output [4:0] out32;
  output [4:0] out33;
  output [4:0] out34;
  output [4:0] out35;
  output [4:0] out36;
  output [4:0] out37;
  output [4:0] out38;
  output [4:0] out39;
  output [4:0] out40;
  output [4:0] out41;
  output [4:0] out42;
  output [4:0] out43;
  output [4:0] out44;
  output [4:0] out45;
  output [4:0] out46;
  output [4:0] out47;
  output [9:0] count2;
  input [4:0] in;
  input reset, clk, test_si, test_se;
  output count1;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n504, n505, n594, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263;
  wire   [9:0] count;

  SIPO_DW01_inc_0 add_143 ( .A(count2), .SUM({N24, N23, N22, N21, N20, N19, 
        N18, N17, N16, N15}) );
  SIPO_DW01_inc_1 add_140 ( .A(count), .SUM({N13, N12, N11, N10, N9, N8, N7, 
        N6, N5, N4}) );
  SDFFRQXLTH count_reg_9_ ( .D(n487), .SI(n1555), .SE(n1497), .CK(clk), .RN(
        n685), .Q(count[9]) );
  SDFFRQXLTH count_reg_8_ ( .D(n486), .SI(count[7]), .SE(n1498), .CK(clk), 
        .RN(n684), .Q(count[8]) );
  SDFFRQXLTH out47_reg_2_ ( .D(n334), .SI(n1553), .SE(n1506), .CK(clk), .RN(
        n679), .Q(out47[2]) );
  SDFFRQXLTH out0_reg_2_ ( .D(n381), .SI(n2257), .SE(n1506), .CK(clk), .RN(
        n675), .Q(out0[2]) );
  SDFFRQXLTH out1_reg_2_ ( .D(n380), .SI(n2011), .SE(n1496), .CK(clk), .RN(
        n675), .Q(out1[2]) );
  SDFFRQXLTH out2_reg_2_ ( .D(n379), .SI(n2128), .SE(n1496), .CK(clk), .RN(
        n675), .Q(out2[2]) );
  SDFFRQXLTH out3_reg_2_ ( .D(n378), .SI(n2014), .SE(n1495), .CK(clk), .RN(
        n675), .Q(out3[2]) );
  SDFFRQXLTH out4_reg_2_ ( .D(n377), .SI(n2017), .SE(n1494), .CK(clk), .RN(
        n675), .Q(out4[2]) );
  SDFFRQXLTH out5_reg_2_ ( .D(n376), .SI(n2242), .SE(n1493), .CK(clk), .RN(
        n675), .Q(out5[2]) );
  SDFFRQXLTH out6_reg_2_ ( .D(n375), .SI(n2137), .SE(n1492), .CK(clk), .RN(
        n675), .Q(out6[2]) );
  SDFFRQXLTH out7_reg_2_ ( .D(n374), .SI(n2020), .SE(n1491), .CK(clk), .RN(
        n675), .Q(out7[2]) );
  SDFFRQXLTH out8_reg_2_ ( .D(n373), .SI(n2023), .SE(n1472), .CK(clk), .RN(
        n675), .Q(out8[2]) );
  SDFFRQXLTH out9_reg_2_ ( .D(n372), .SI(n2230), .SE(n1471), .CK(clk), .RN(
        n680), .Q(out9[2]) );
  SDFFRQXLTH out10_reg_2_ ( .D(n371), .SI(n2233), .SE(n1470), .CK(clk), .RN(
        n692), .Q(out10[2]) );
  SDFFRQXLTH out11_reg_2_ ( .D(n370), .SI(n2146), .SE(n1469), .CK(clk), .RN(
        n691), .Q(out11[2]) );
  SDFFRQXLTH out13_reg_2_ ( .D(n368), .SI(n2029), .SE(n1467), .CK(clk), .RN(
        n691), .Q(out13[2]) );
  SDFFRQXLTH out15_reg_2_ ( .D(n366), .SI(n2035), .SE(n1466), .CK(clk), .RN(
        n691), .Q(out15[2]) );
  SDFFRQXLTH out16_reg_2_ ( .D(n365), .SI(n2101), .SE(n1467), .CK(clk), .RN(
        n691), .Q(out16[2]) );
  SDFFRQXLTH out17_reg_2_ ( .D(n364), .SI(n2038), .SE(n1478), .CK(clk), .RN(
        n691), .Q(out17[2]) );
  SDFFRQXLTH out18_reg_2_ ( .D(n363), .SI(n2041), .SE(n1477), .CK(clk), .RN(
        n691), .Q(out18[2]) );
  SDFFRQXLTH out19_reg_2_ ( .D(n362), .SI(n2044), .SE(n1476), .CK(clk), .RN(
        n691), .Q(out19[2]) );
  SDFFRQXLTH out20_reg_2_ ( .D(n361), .SI(n2047), .SE(n1475), .CK(clk), .RN(
        n691), .Q(out20[2]) );
  SDFFRQXLTH out21_reg_2_ ( .D(n360), .SI(n2104), .SE(n1474), .CK(clk), .RN(
        n691), .Q(out21[2]) );
  SDFFRQXLTH out22_reg_2_ ( .D(n359), .SI(n2050), .SE(n1549), .CK(clk), .RN(
        n691), .Q(out22[2]) );
  SDFFRQXLTH out23_reg_2_ ( .D(n358), .SI(n2131), .SE(n1549), .CK(clk), .RN(
        n691), .Q(out23[2]) );
  SDFFRQXLTH out24_reg_2_ ( .D(n357), .SI(n2053), .SE(n1549), .CK(clk), .RN(
        n690), .Q(out24[2]) );
  SDFFRQXLTH out25_reg_2_ ( .D(n356), .SI(n2245), .SE(n1466), .CK(clk), .RN(
        n690), .Q(out25[2]) );
  SDFFRQXLTH out27_reg_2_ ( .D(n354), .SI(n2056), .SE(n1484), .CK(clk), .RN(
        n690), .Q(out27[2]) );
  SDFFRQXLTH out29_reg_2_ ( .D(n352), .SI(n2062), .SE(n1482), .CK(clk), .RN(
        n690), .Q(out29[2]) );
  SDFFRQXLTH out30_reg_2_ ( .D(n351), .SI(n2065), .SE(n1481), .CK(clk), .RN(
        n690), .Q(out30[2]) );
  SDFFRQXLTH out31_reg_2_ ( .D(n350), .SI(n2227), .SE(n1480), .CK(clk), .RN(
        n690), .Q(out31[2]) );
  SDFFRQXLTH out33_reg_2_ ( .D(n348), .SI(n2071), .SE(n1550), .CK(clk), .RN(
        n690), .Q(out33[2]) );
  SDFFRQXLTH out34_reg_2_ ( .D(n347), .SI(n2134), .SE(n1550), .CK(clk), .RN(
        n690), .Q(out34[2]) );
  SDFFRQXLTH out35_reg_2_ ( .D(n346), .SI(n2074), .SE(n1467), .CK(clk), .RN(
        n690), .Q(out35[2]) );
  SDFFRQXLTH out36_reg_2_ ( .D(n345), .SI(n2077), .SE(n1467), .CK(clk), .RN(
        n690), .Q(out36[2]) );
  SDFFRQXLTH out37_reg_2_ ( .D(n344), .SI(n2236), .SE(n1490), .CK(clk), .RN(
        n690), .Q(out37[2]) );
  SDFFRQXLTH out38_reg_2_ ( .D(n343), .SI(n2140), .SE(n1489), .CK(clk), .RN(
        n689), .Q(out38[2]) );
  SDFFRQXLTH out39_reg_2_ ( .D(n342), .SI(n2080), .SE(n1488), .CK(clk), .RN(
        n689), .Q(out39[2]) );
  SDFFRQXLTH out40_reg_2_ ( .D(n341), .SI(n2239), .SE(n1487), .CK(clk), .RN(
        n689), .Q(out40[2]) );
  SDFFRQXLTH out41_reg_2_ ( .D(n340), .SI(n2125), .SE(n1486), .CK(clk), .RN(
        n689), .Q(out41[2]) );
  SDFFRQXLTH out42_reg_2_ ( .D(n339), .SI(n2083), .SE(n1551), .CK(clk), .RN(
        n689), .Q(out42[2]) );
  SDFFRQXLTH out43_reg_2_ ( .D(n338), .SI(n2221), .SE(n1551), .CK(clk), .RN(
        n689), .Q(out43[2]) );
  SDFFRQXLTH out44_reg_2_ ( .D(n337), .SI(n2224), .SE(n1551), .CK(clk), .RN(
        n689), .Q(out44[2]) );
  SDFFRQXLTH out46_reg_2_ ( .D(n335), .SI(n1573), .SE(n1506), .CK(clk), .RN(
        n689), .Q(out46[2]) );
  SDFFRQXLTH out26_reg_2_ ( .D(n355), .SI(n2143), .SE(n1466), .CK(clk), .RN(
        n685), .Q(out26[2]) );
  SDFFRQX2TH out26_reg_0_ ( .D(n259), .SI(n2209), .SE(n1500), .CK(clk), .RN(
        n677), .Q(out26[0]) );
  SDFFRQXLTH out12_reg_2_ ( .D(n369), .SI(n2026), .SE(n1466), .CK(clk), .RN(
        n691), .Q(out12[2]) );
  SDFFRQXLTH out14_reg_2_ ( .D(n367), .SI(n2032), .SE(n1499), .CK(clk), .RN(
        n691), .Q(out14[2]) );
  SDFFRQXLTH out28_reg_2_ ( .D(n353), .SI(n2059), .SE(n1483), .CK(clk), .RN(
        n690), .Q(out28[2]) );
  SDFFRQX1TH out4_reg_4_ ( .D(n473), .SI(n1849), .SE(n1471), .CK(clk), .RN(
        n677), .Q(out4[4]) );
  SDFFRQX1TH out8_reg_4_ ( .D(n469), .SI(n1948), .SE(n1473), .CK(clk), .RN(
        n676), .Q(out8[4]) );
  SDFFRQX1TH out32_reg_4_ ( .D(n445), .SI(n1963), .SE(n1540), .CK(clk), .RN(
        n686), .Q(out32[4]) );
  SDFFRQX1TH out19_reg_4_ ( .D(n458), .SI(n1855), .SE(n1532), .CK(clk), .RN(
        n687), .Q(out19[4]) );
  SDFFRQX1TH out13_reg_4_ ( .D(n464), .SI(n1840), .SE(n1476), .CK(clk), .RN(
        n679), .Q(out13[4]) );
  SDFFRQX1TH out1_reg_4_ ( .D(n476), .SI(n1945), .SE(n1469), .CK(clk), .RN(
        n688), .Q(out1[4]) );
  SDFFRQX1TH out20_reg_4_ ( .D(n457), .SI(n1858), .SE(n1533), .CK(clk), .RN(
        n687), .Q(out20[4]) );
  SDFFRQX1TH out12_reg_4_ ( .D(n465), .SI(n1969), .SE(n1528), .CK(clk), .RN(
        n683), .Q(out12[4]) );
  SDFFRQX1TH out36_reg_4_ ( .D(n441), .SI(n1867), .SE(n1490), .CK(clk), .RN(
        n686), .Q(out36[4]) );
  SDFFRQX1TH out28_reg_4_ ( .D(n449), .SI(n1864), .SE(n1485), .CK(clk), .RN(
        n687), .Q(out28[4]) );
  SDFFRQX1TH out14_reg_4_ ( .D(n463), .SI(n1843), .SE(n1529), .CK(clk), .RN(
        n691), .Q(out14[4]) );
  SDFFRQX1TH out30_reg_1_ ( .D(n303), .SI(n1660), .SE(n1486), .CK(clk), .RN(
        n693), .Q(out30[1]) );
  SDFFRQX1TH out3_reg_1_ ( .D(n330), .SI(n1588), .SE(n1470), .CK(clk), .RN(
        n689), .Q(out3[1]) );
  SDFFRQX1TH out15_reg_1_ ( .D(n318), .SI(n1624), .SE(n1477), .CK(clk), .RN(
        n701), .Q(out15[1]) );
  SDFFRQX1TH out22_reg_1_ ( .D(n311), .SI(n1642), .SE(n1481), .CK(clk), .RN(
        n694), .Q(out22[1]) );
  SDFFRQX1TH out24_reg_1_ ( .D(n309), .SI(n1645), .SE(n1535), .CK(clk), .RN(
        n695), .Q(out24[1]) );
  SDFFRQX1TH out17_reg_1_ ( .D(n316), .SI(n1627), .SE(n1478), .CK(clk), .RN(
        n675), .Q(out17[1]) );
  SDFFRQX1TH out29_reg_1_ ( .D(n304), .SI(n1657), .SE(n1538), .CK(clk), .RN(
        n699), .Q(out29[1]) );
  SDFFRQX1TH out46_reg_1_ ( .D(n287), .SI(n1564), .SE(n1548), .CK(clk), .RN(
        n688), .Q(out46[1]) );
  SDFFRQX1TH out18_reg_1_ ( .D(n315), .SI(n1630), .SE(n1531), .CK(clk), .RN(
        n698), .Q(out18[1]) );
  SDFFRQX1TH out35_reg_1_ ( .D(n298), .SI(n1672), .SE(n1489), .CK(clk), .RN(
        n688), .Q(out35[1]) );
  SDFFRQX1TH out7_reg_1_ ( .D(n326), .SI(n1609), .SE(n1525), .CK(clk), .RN(
        n685), .Q(out7[1]) );
  SDFFRQX1TH out33_reg_1_ ( .D(n300), .SI(n1669), .SE(n1540), .CK(clk), .RN(
        n699), .Q(out33[1]) );
  SDFFRQX1TH out39_reg_1_ ( .D(n294), .SI(n1681), .SE(n1544), .CK(clk), .RN(
        n688), .Q(out39[1]) );
  SDFFRQX1TH out8_reg_1_ ( .D(n325), .SI(n1612), .SE(n1525), .CK(clk), .RN(
        reset), .Q(out8[1]) );
  SDFFRQX1TH out27_reg_1_ ( .D(n306), .SI(n1651), .SE(n1484), .CK(clk), .RN(
        n700), .Q(out27[1]) );
  SDFFRQX1TH out4_reg_1_ ( .D(n329), .SI(n1600), .SE(n1523), .CK(clk), .RN(
        n689), .Q(out4[1]) );
  SDFFRQX1TH out19_reg_1_ ( .D(n314), .SI(n1633), .SE(n1532), .CK(clk), .RN(
        n697), .Q(out19[1]) );
  SDFFRQX1TH out13_reg_1_ ( .D(n320), .SI(n1618), .SE(n1528), .CK(clk), .RN(
        n700), .Q(out13[1]) );
  SDFFRQX1TH out12_reg_1_ ( .D(n321), .SI(n1615), .SE(n1475), .CK(clk), .RN(
        n703), .Q(out12[1]) );
  SDFFRQX1TH out20_reg_1_ ( .D(n313), .SI(n1636), .SE(n1480), .CK(clk), .RN(
        n685), .Q(out20[1]) );
  SDFFRQX1TH out1_reg_1_ ( .D(n332), .SI(n1597), .SE(n1521), .CK(clk), .RN(
        n689), .Q(out1[1]) );
  SDFFRQX1TH out36_reg_1_ ( .D(n297), .SI(n1675), .SE(n1542), .CK(clk), .RN(
        n688), .Q(out36[1]) );
  SDFFRQX1TH out28_reg_1_ ( .D(n305), .SI(n1654), .SE(n1537), .CK(clk), .RN(
        n698), .Q(out28[1]) );
  SDFFRQX2TH out3_reg_0_ ( .D(n282), .SI(n2206), .SE(n1511), .CK(clk), .RN(
        n679), .Q(out3[0]) );
  SDFFRQX2TH out21_reg_0_ ( .D(n264), .SI(n1999), .SE(n1499), .CK(clk), .RN(
        n677), .Q(out21[0]) );
  SDFFRQX2TH out6_reg_0_ ( .D(n279), .SI(n2212), .SE(n1509), .CK(clk), .RN(
        n678), .Q(out6[0]) );
  SDFFRQX2TH out44_reg_0_ ( .D(n241), .SI(n2170), .SE(n1504), .CK(clk), .RN(
        n676), .Q(out44[0]) );
  SDFFRQX2TH out31_reg_0_ ( .D(n254), .SI(n2203), .SE(n1501), .CK(clk), .RN(
        n677), .Q(out31[0]) );
  SDFFRQX2TH out38_reg_0_ ( .D(n247), .SI(n2158), .SE(n1518), .CK(clk), .RN(
        n676), .Q(out38[0]) );
  SDFFRQX2TH out25_reg_0_ ( .D(n260), .SI(n2164), .SE(n1500), .CK(clk), .RN(
        n677), .Q(out25[0]) );
  SDFFRQX2TH out0_reg_0_ ( .D(n285), .SI(n1558), .SE(n1511), .CK(clk), .RN(
        n679), .Q(out0[0]) );
  SDFFRQX2TH out40_reg_0_ ( .D(n245), .SI(n2095), .SE(n1503), .CK(clk), .RN(
        n676), .Q(out40[0]) );
  SDFFRQX2TH out5_reg_0_ ( .D(n280), .SI(n1981), .SE(n1509), .CK(clk), .RN(
        n678), .Q(out5[0]) );
  SDFFRQX2TH out43_reg_0_ ( .D(n242), .SI(n2167), .SE(n1519), .CK(clk), .RN(
        n676), .Q(out43[0]) );
  SDFFRQX2TH out42_reg_0_ ( .D(n243), .SI(n2176), .SE(n1519), .CK(clk), .RN(
        n676), .Q(out42[0]) );
  SDFFRQX2TH out30_reg_0_ ( .D(n255), .SI(n2155), .SE(n1501), .CK(clk), .RN(
        n677), .Q(out30[0]) );
  SDFFRQX2TH out22_reg_0_ ( .D(n263), .SI(n2188), .SE(n1515), .CK(clk), .RN(
        n677), .Q(out22[0]) );
  SDFFRQX2TH out15_reg_0_ ( .D(n270), .SI(n1993), .SE(n1498), .CK(clk), .RN(
        n678), .Q(out15[0]) );
  SDFFRQX2TH out24_reg_0_ ( .D(n261), .SI(n2161), .SE(n1515), .CK(clk), .RN(
        n677), .Q(out24[0]) );
  SDFFRQX2TH out17_reg_0_ ( .D(n268), .SI(n2089), .SE(n1514), .CK(clk), .RN(
        n701), .Q(out17[0]) );
  SDFFRQX2TH out29_reg_0_ ( .D(n256), .SI(n2002), .SE(n1516), .CK(clk), .RN(
        n677), .Q(out29[0]) );
  SDFFRQX2TH out46_reg_0_ ( .D(n239), .SI(n2098), .SE(n1520), .CK(clk), .RN(
        n679), .Q(out46[0]) );
  SDFFRQX2TH out18_reg_0_ ( .D(n267), .SI(n2152), .SE(n1514), .CK(clk), .RN(
        n678), .Q(out18[0]) );
  SDFFRQX2TH out7_reg_0_ ( .D(n278), .SI(n2218), .SE(n1512), .CK(clk), .RN(
        n678), .Q(out7[0]) );
  SDFFRQX2TH out35_reg_0_ ( .D(n250), .SI(n2185), .SE(n1502), .CK(clk), .RN(
        n676), .Q(out35[0]) );
  SDFFRQX2TH out39_reg_0_ ( .D(n246), .SI(n2215), .SE(n1518), .CK(clk), .RN(
        n676), .Q(out39[0]) );
  SDFFRQX2TH out8_reg_0_ ( .D(n277), .SI(n1978), .SE(n1512), .CK(clk), .RN(
        n678), .Q(out8[0]) );
  SDFFRQX2TH out33_reg_0_ ( .D(n252), .SI(n2005), .SE(n1517), .CK(clk), .RN(
        n676), .Q(out33[0]) );
  SDFFRQX2TH out27_reg_0_ ( .D(n258), .SI(n2194), .SE(n1516), .CK(clk), .RN(
        n677), .Q(out27[0]) );
  SDFFRQX2TH out19_reg_0_ ( .D(n266), .SI(n2116), .SE(n1514), .CK(clk), .RN(
        n677), .Q(out19[0]) );
  SDFFRQX2TH out4_reg_0_ ( .D(n281), .SI(n2110), .SE(n1509), .CK(clk), .RN(
        n679), .Q(out4[0]) );
  SDFFRQX2TH out12_reg_0_ ( .D(n273), .SI(n2119), .SE(n1513), .CK(clk), .RN(
        n678), .Q(out12[0]) );
  SDFFRQX2TH out20_reg_0_ ( .D(n265), .SI(n1996), .SE(n1499), .CK(clk), .RN(
        n685), .Q(out20[0]) );
  SDFFRQX2TH out28_reg_0_ ( .D(n257), .SI(n2092), .SE(n1516), .CK(clk), .RN(
        n677), .Q(out28[0]) );
  SDFFRQX1TH out14_reg_1_ ( .D(n319), .SI(n1621), .SE(n1529), .CK(clk), .RN(
        n692), .Q(out14[1]) );
  SDFFRQX2TH out1_reg_0_ ( .D(n284), .SI(n2263), .SE(n1511), .CK(clk), .RN(
        n679), .Q(out1[0]) );
  SDFFRQX2TH out13_reg_0_ ( .D(n272), .SI(n1987), .SE(n1513), .CK(clk), .RN(
        n678), .Q(out13[0]) );
  SDFFRQX2TH out14_reg_0_ ( .D(n271), .SI(n1990), .SE(n1513), .CK(clk), .RN(
        n678), .Q(out14[0]) );
  SDFFRQX2TH out36_reg_0_ ( .D(n249), .SI(n2122), .SE(n1502), .CK(clk), .RN(
        n676), .Q(out36[0]) );
  SDFFRQX1TH count_reg_1_ ( .D(n479), .SI(n1552), .SE(n1468), .CK(clk), .RN(
        n684), .Q(count[1]) );
  SDFFRQX1TH count_reg_2_ ( .D(n480), .SI(count[1]), .SE(n1468), .CK(clk), 
        .RN(n684), .Q(count[2]) );
  SDFFRQX1TH count_reg_3_ ( .D(n481), .SI(count[2]), .SE(test_se), .CK(clk), 
        .RN(n684), .Q(count[3]) );
  SDFFRQX1TH count_reg_4_ ( .D(n482), .SI(count[3]), .SE(n1504), .CK(clk), 
        .RN(n684), .Q(count[4]) );
  SDFFRQX1TH count_reg_5_ ( .D(n483), .SI(count[4]), .SE(n1503), .CK(clk), 
        .RN(n684), .Q(count[5]) );
  SDFFRQX1TH count_reg_6_ ( .D(n484), .SI(count[5]), .SE(n1502), .CK(clk), 
        .RN(n684), .Q(count[6]) );
  SDFFRQX1TH count_reg_0_ ( .D(n488), .SI(count2[9]), .SE(n1520), .CK(clk), 
        .RN(n684), .Q(count[0]) );
  SDFFRQX1TH out14_reg_3_ ( .D(n415), .SI(n1582), .SE(n1529), .CK(clk), .RN(
        n682), .Q(out14[3]) );
  SDFFRQX1TH out4_reg_3_ ( .D(n425), .SI(n1708), .SE(n1523), .CK(clk), .RN(
        n683), .Q(out4[3]) );
  SDFFRQX1TH out19_reg_3_ ( .D(n410), .SI(n1747), .SE(n1532), .CK(clk), .RN(
        n681), .Q(out19[3]) );
  SDFFRQX1TH out20_reg_3_ ( .D(n409), .SI(n1750), .SE(n1480), .CK(clk), .RN(
        n681), .Q(out20[3]) );
  SDFFRQX1TH out28_reg_3_ ( .D(n401), .SI(n1585), .SE(n1485), .CK(clk), .RN(
        n681), .Q(out28[3]) );
  SDFFRQX1TH out36_reg_3_ ( .D(n393), .SI(n1792), .SE(n1542), .CK(clk), .RN(
        n680), .Q(out36[3]) );
  SDFFRQX1TH out3_reg_3_ ( .D(n426), .SI(n1705), .SE(n1470), .CK(clk), .RN(
        n683), .Q(out3[3]) );
  SDFFRQX1TH out5_reg_3_ ( .D(n424), .SI(n1711), .SE(n1524), .CK(clk), .RN(
        n683), .Q(out5[3]) );
  SDFFRQX1TH out6_reg_3_ ( .D(n423), .SI(n1714), .SE(n1472), .CK(clk), .RN(
        n682), .Q(out6[3]) );
  SDFFRQX1TH out7_reg_3_ ( .D(n422), .SI(n1717), .SE(n1525), .CK(clk), .RN(
        n682), .Q(out7[3]) );
  SDFFRQX1TH out15_reg_3_ ( .D(n414), .SI(n1735), .SE(n1477), .CK(clk), .RN(
        n682), .Q(out15[3]) );
  SDFFRQX1TH out21_reg_3_ ( .D(n408), .SI(n1753), .SE(n1533), .CK(clk), .RN(
        n681), .Q(out21[3]) );
  SDFFRQX1TH out22_reg_3_ ( .D(n407), .SI(n1756), .SE(n1534), .CK(clk), .RN(
        n681), .Q(out22[3]) );
  SDFFRQX1TH out24_reg_3_ ( .D(n405), .SI(n1762), .SE(n1535), .CK(clk), .RN(
        n681), .Q(out24[3]) );
  SDFFRQX1TH out25_reg_3_ ( .D(n404), .SI(n1765), .SE(n1483), .CK(clk), .RN(
        n681), .Q(out25[3]) );
  SDFFRQX1TH out26_reg_3_ ( .D(n403), .SI(n1768), .SE(n1536), .CK(clk), .RN(
        n681), .Q(out26[3]) );
  SDFFRQX1TH out30_reg_3_ ( .D(n399), .SI(n1777), .SE(n1486), .CK(clk), .RN(
        n681), .Q(out30[3]) );
  SDFFRQX1TH out31_reg_3_ ( .D(n398), .SI(n1780), .SE(n1539), .CK(clk), .RN(
        n681), .Q(out31[3]) );
  SDFFRQX1TH out35_reg_3_ ( .D(n394), .SI(n1789), .SE(n1489), .CK(clk), .RN(
        n680), .Q(out35[3]) );
  SDFFRQX1TH out38_reg_3_ ( .D(n391), .SI(n1798), .SE(n1491), .CK(clk), .RN(
        n680), .Q(out38[3]) );
  SDFFRQX1TH out39_reg_3_ ( .D(n390), .SI(n1801), .SE(n1544), .CK(clk), .RN(
        n680), .Q(out39[3]) );
  SDFFRQX1TH out40_reg_3_ ( .D(n389), .SI(n1804), .SE(n1492), .CK(clk), .RN(
        n680), .Q(out40[3]) );
  SDFFRQX1TH out42_reg_3_ ( .D(n387), .SI(n1810), .SE(n1493), .CK(clk), .RN(
        n680), .Q(out42[3]) );
  SDFFRQX1TH out43_reg_3_ ( .D(n386), .SI(n1813), .SE(n1546), .CK(clk), .RN(
        n680), .Q(out43[3]) );
  SDFFRQX1TH out44_reg_3_ ( .D(n385), .SI(n1816), .SE(n1547), .CK(clk), .RN(
        n679), .Q(out44[3]) );
  SDFFRQX1TH out46_reg_3_ ( .D(n383), .SI(n1567), .SE(n1548), .CK(clk), .RN(
        n679), .Q(out46[3]) );
  SDFFRQX1TH out2_reg_3_ ( .D(n427), .SI(n1702), .SE(n1522), .CK(clk), .RN(
        n683), .Q(out2[3]) );
  SDFFRQX1TH out10_reg_3_ ( .D(n419), .SI(n1726), .SE(n1474), .CK(clk), .RN(
        n682), .Q(out10[3]) );
  SDFFRQX1TH out11_reg_3_ ( .D(n418), .SI(n1729), .SE(n1527), .CK(clk), .RN(
        n682), .Q(out11[3]) );
  SDFFRQX1TH out17_reg_3_ ( .D(n412), .SI(n1741), .SE(n1531), .CK(clk), .RN(
        n682), .Q(out17[3]) );
  SDFFRQX1TH out23_reg_3_ ( .D(n406), .SI(n1759), .SE(n1482), .CK(clk), .RN(
        n681), .Q(out23[3]) );
  SDFFRQX1TH out29_reg_3_ ( .D(n400), .SI(n1774), .SE(n1538), .CK(clk), .RN(
        n681), .Q(out29[3]) );
  SDFFRQX1TH out33_reg_3_ ( .D(n396), .SI(n1783), .SE(n1488), .CK(clk), .RN(
        n680), .Q(out33[3]) );
  SDFFRQX1TH out37_reg_3_ ( .D(n392), .SI(n1795), .SE(n1543), .CK(clk), .RN(
        n680), .Q(out37[3]) );
  SDFFRQX1TH out41_reg_3_ ( .D(n388), .SI(n1807), .SE(n1545), .CK(clk), .RN(
        n680), .Q(out41[3]) );
  SDFFRQXLTH out45_reg_2_ ( .D(n336), .SI(n2107), .SE(n1506), .CK(clk), .RN(
        n689), .Q(out45[2]) );
  SDFFRQXLTH out32_reg_2_ ( .D(n349), .SI(n2068), .SE(n1550), .CK(clk), .RN(
        n690), .Q(out32[2]) );
  SDFFRQX1TH out8_reg_3_ ( .D(n421), .SI(n1720), .SE(n1473), .CK(clk), .RN(
        n682), .Q(out8[3]) );
  SDFFRQX1TH out13_reg_3_ ( .D(n416), .SI(n1732), .SE(n1476), .CK(clk), .RN(
        n682), .Q(out13[3]) );
  SDFFRQX1TH out32_reg_3_ ( .D(n397), .SI(n1690), .SE(n1540), .CK(clk), .RN(
        n680), .Q(out32[3]) );
  SDFFRQX1TH out1_reg_3_ ( .D(n428), .SI(n1699), .SE(n1469), .CK(clk), .RN(
        n683), .Q(out1[3]) );
  SDFFRQX1TH out27_reg_3_ ( .D(n402), .SI(n1771), .SE(n1537), .CK(clk), .RN(
        n681), .Q(out27[3]) );
  SDFFRQX1TH out0_reg_3_ ( .D(n429), .SI(n2251), .SE(n1521), .CK(clk), .RN(
        n683), .Q(out0[3]) );
  SDFFRQX1TH out12_reg_3_ ( .D(n417), .SI(n1579), .SE(n1528), .CK(clk), .RN(
        n682), .Q(out12[3]) );
  SDFFRQX1TH out16_reg_3_ ( .D(n413), .SI(n1738), .SE(n1530), .CK(clk), .RN(
        n682), .Q(out16[3]) );
  SDFFRQX1TH out45_reg_3_ ( .D(n384), .SI(n1693), .SE(n1495), .CK(clk), .RN(
        n679), .Q(out45[3]) );
  SDFFRQX1TH out11_reg_4_ ( .D(n466), .SI(n1957), .SE(n1475), .CK(clk), .RN(
        n690), .Q(out11[4]) );
  SDFFRQX1TH out18_reg_4_ ( .D(n459), .SI(n1852), .SE(n1479), .CK(clk), .RN(
        n687), .Q(out18[4]) );
  SDFFRQX1TH out29_reg_4_ ( .D(n448), .SI(n1909), .SE(n1538), .CK(clk), .RN(
        n687), .Q(out29[4]) );
  SDFFRQX1TH out37_reg_4_ ( .D(n440), .SI(n1918), .SE(n1543), .CK(clk), .RN(
        n686), .Q(out37[4]) );
  SDFFRQX1TH out24_reg_4_ ( .D(n453), .SI(n1894), .SE(n1535), .CK(clk), .RN(
        n687), .Q(out24[4]) );
  SDFFRQX1TH out43_reg_4_ ( .D(n434), .SI(n1936), .SE(n1494), .CK(clk), .RN(
        n686), .Q(out43[4]) );
  SDFFRQX1TH out41_reg_4_ ( .D(n436), .SI(n1930), .SE(n1493), .CK(clk), .RN(
        n686), .Q(out41[4]) );
  SDFFRQX1TH out40_reg_4_ ( .D(n437), .SI(n1927), .SE(n1545), .CK(clk), .RN(
        n686), .Q(out40[4]) );
  SDFFRQX1TH out42_reg_4_ ( .D(n435), .SI(n1933), .SE(n1546), .CK(clk), .RN(
        n686), .Q(out42[4]) );
  SDFFRQX1TH out9_reg_4_ ( .D(n468), .SI(n1951), .SE(n1526), .CK(clk), .RN(
        n689), .Q(out9[4]) );
  SDFFRQX1TH out46_reg_4_ ( .D(n431), .SI(n1570), .SE(n1548), .CK(clk), .RN(
        n685), .Q(out46[4]) );
  SDFFRQX1TH out15_reg_4_ ( .D(n462), .SI(n1882), .SE(n1530), .CK(clk), .RN(
        n680), .Q(out15[4]) );
  SDFFRQX1TH out35_reg_4_ ( .D(n442), .SI(n1870), .SE(n1542), .CK(clk), .RN(
        n686), .Q(out35[4]) );
  SDFFRQX1TH out21_reg_4_ ( .D(n456), .SI(n1888), .SE(n1481), .CK(clk), .RN(
        n687), .Q(out21[4]) );
  SDFFRQX1TH out44_reg_4_ ( .D(n433), .SI(n1939), .SE(n1547), .CK(clk), .RN(
        n685), .Q(out44[4]) );
  SDFFRQX1TH out27_reg_4_ ( .D(n450), .SI(n1861), .SE(n1537), .CK(clk), .RN(
        n687), .Q(out27[4]) );
  SDFFRQX1TH out22_reg_4_ ( .D(n455), .SI(n1891), .SE(n1534), .CK(clk), .RN(
        n687), .Q(out22[4]) );
  SDFFRQX1TH out17_reg_4_ ( .D(n460), .SI(n1885), .SE(n1531), .CK(clk), .RN(
        n685), .Q(out17[4]) );
  SDFFRQX1TH out33_reg_4_ ( .D(n444), .SI(n1966), .SE(n1488), .CK(clk), .RN(
        n686), .Q(out33[4]) );
  SDFFRQX1TH out30_reg_4_ ( .D(n447), .SI(n1906), .SE(n1539), .CK(clk), .RN(
        n687), .Q(out30[4]) );
  SDFFRQX1TH out23_reg_4_ ( .D(n454), .SI(n1897), .SE(n1482), .CK(clk), .RN(
        n687), .Q(out23[4]) );
  SDFFRQX1TH out10_reg_4_ ( .D(n467), .SI(n1954), .SE(n1527), .CK(clk), .RN(
        n688), .Q(out10[4]) );
  SDFFRQX1TH out2_reg_4_ ( .D(n475), .SI(n1873), .SE(n1522), .CK(clk), .RN(
        n688), .Q(out2[4]) );
  SDFFRQX1TH out25_reg_4_ ( .D(n452), .SI(n1900), .SE(n1536), .CK(clk), .RN(
        n687), .Q(out25[4]) );
  SDFFRQX1TH out5_reg_4_ ( .D(n472), .SI(n1876), .SE(n1524), .CK(clk), .RN(
        n686), .Q(out5[4]) );
  SDFFRQX1TH out39_reg_4_ ( .D(n438), .SI(n1924), .SE(n1544), .CK(clk), .RN(
        n686), .Q(out39[4]) );
  SDFFRQX1TH out34_reg_4_ ( .D(n443), .SI(n1915), .SE(n1541), .CK(clk), .RN(
        n686), .Q(out34[4]) );
  SDFFRQX1TH out26_reg_4_ ( .D(n451), .SI(n1903), .SE(n1484), .CK(clk), .RN(
        n687), .Q(out26[4]) );
  SDFFRQX1TH out6_reg_4_ ( .D(n471), .SI(n1879), .SE(n1472), .CK(clk), .RN(
        n687), .Q(out6[4]) );
  SDFFRQX1TH out3_reg_4_ ( .D(n474), .SI(n1846), .SE(n1523), .CK(clk), .RN(
        n694), .Q(out3[4]) );
  SDFFRQX1TH out38_reg_4_ ( .D(n439), .SI(n1921), .SE(n1491), .CK(clk), .RN(
        n686), .Q(out38[4]) );
  SDFFRQX1TH out16_reg_4_ ( .D(n461), .SI(n1960), .SE(n1478), .CK(clk), .RN(
        n694), .Q(out16[4]) );
  SDFFRQX1TH out31_reg_4_ ( .D(n446), .SI(n1912), .SE(n1487), .CK(clk), .RN(
        n686), .Q(out31[4]) );
  SDFFRQX1TH out47_reg_4_ ( .D(n430), .SI(out47[3]), .SE(n1468), .CK(clk), 
        .RN(n675), .Q(out47[4]) );
  SDFFRQX1TH out44_reg_1_ ( .D(n289), .SI(n1591), .SE(n1494), .CK(clk), .RN(
        n685), .Q(out44[1]) );
  SDFFRQX1TH out31_reg_1_ ( .D(n302), .SI(n1663), .SE(n1539), .CK(clk), .RN(
        n697), .Q(out31[1]) );
  SDFFRQX1TH out2_reg_1_ ( .D(n331), .SI(n1822), .SE(n1522), .CK(clk), .RN(
        n689), .Q(out2[1]) );
  SDFFRQX1TH out9_reg_1_ ( .D(n324), .SI(n1972), .SE(n1526), .CK(clk), .RN(
        n702), .Q(out9[1]) );
  SDFFRQX1TH out10_reg_1_ ( .D(n323), .SI(n1975), .SE(n1474), .CK(clk), .RN(
        n695), .Q(out10[1]) );
  SDFFRQX1TH out23_reg_1_ ( .D(n310), .SI(n1831), .SE(n1534), .CK(clk), .RN(
        n696), .Q(out23[1]) );
  SDFFRQX1TH out34_reg_1_ ( .D(n299), .SI(n1834), .SE(n1541), .CK(clk), .RN(
        n688), .Q(out34[1]) );
  SDFFRQX1TH out37_reg_1_ ( .D(n296), .SI(n1825), .SE(n1490), .CK(clk), .RN(
        n688), .Q(out37[1]) );
  SDFFRQX1TH out41_reg_1_ ( .D(n292), .SI(n1828), .SE(n1545), .CK(clk), .RN(
        n688), .Q(out41[1]) );
  SDFFRQX1TH out43_reg_1_ ( .D(n290), .SI(n1687), .SE(n1546), .CK(clk), .RN(
        n688), .Q(out43[1]) );
  SDFFRQX1TH out40_reg_1_ ( .D(n293), .SI(n1684), .SE(n1492), .CK(clk), .RN(
        n688), .Q(out40[1]) );
  SDFFRQX1TH out5_reg_1_ ( .D(n328), .SI(n1603), .SE(n1471), .CK(clk), .RN(
        n704), .Q(out5[1]) );
  SDFFRQX1TH out6_reg_1_ ( .D(n327), .SI(n1606), .SE(n1524), .CK(clk), .RN(
        n674), .Q(out6[1]) );
  SDFFRQX1TH out38_reg_1_ ( .D(n295), .SI(n1678), .SE(n1543), .CK(clk), .RN(
        n685), .Q(out38[1]) );
  SDFFRQX1TH out25_reg_1_ ( .D(n308), .SI(n1648), .SE(n1483), .CK(clk), .RN(
        n704), .Q(out25[1]) );
  SDFFRQX1TH out26_reg_1_ ( .D(n307), .SI(n1819), .SE(n1536), .CK(clk), .RN(
        n674), .Q(out26[1]) );
  SDFFRQX1TH out16_reg_1_ ( .D(n317), .SI(n1696), .SE(n1530), .CK(clk), .RN(
        n693), .Q(out16[1]) );
  SDFFRQX1TH out21_reg_1_ ( .D(n312), .SI(n1639), .SE(n1533), .CK(clk), .RN(
        n696), .Q(out21[1]) );
  SDFFRQX1TH out45_reg_1_ ( .D(n288), .SI(n1594), .SE(n1547), .CK(clk), .RN(
        n688), .Q(out45[1]) );
  SDFFRQX1TH out0_reg_1_ ( .D(n333), .SI(n2248), .SE(n1501), .CK(clk), .RN(
        n675), .Q(out0[1]) );
  SDFFRQX1TH out47_reg_1_ ( .D(n286), .SI(out47[0]), .SE(n1496), .CK(clk), 
        .RN(n676), .Q(out47[1]) );
  SDFFRQX1TH out0_reg_4_ ( .D(n477), .SI(n2254), .SE(n1521), .CK(clk), .RN(
        n679), .Q(out0[4]) );
  SDFFRQX1TH out11_reg_1_ ( .D(n322), .SI(n1837), .SE(n1527), .CK(clk), .RN(
        n685), .Q(out11[1]) );
  SDFFRQX2TH out2_reg_0_ ( .D(n283), .SI(n1561), .SE(n1511), .CK(clk), .RN(
        n679), .Q(out2[0]) );
  SDFFRQX2TH out10_reg_0_ ( .D(n275), .SI(n2179), .SE(n1497), .CK(clk), .RN(
        n678), .Q(out10[0]) );
  SDFFRQX2TH out34_reg_0_ ( .D(n251), .SI(n2200), .SE(n1517), .CK(clk), .RN(
        n676), .Q(out34[0]) );
  SDFFRQX2TH out37_reg_0_ ( .D(n248), .SI(n2008), .SE(n1518), .CK(clk), .RN(
        n676), .Q(out37[0]) );
  SDFFRQX2TH out9_reg_0_ ( .D(n276), .SI(n1984), .SE(n1512), .CK(clk), .RN(
        n678), .Q(out9[0]) );
  SDFFRQX2TH out23_reg_0_ ( .D(n262), .SI(n2197), .SE(n1515), .CK(clk), .RN(
        n677), .Q(out23[0]) );
  SDFFRQX2TH out16_reg_0_ ( .D(n269), .SI(n2182), .SE(n1498), .CK(clk), .RN(
        n678), .Q(out16[0]) );
  SDFFRQX2TH out41_reg_0_ ( .D(n244), .SI(n2173), .SE(n1503), .CK(clk), .RN(
        n676), .Q(out41[0]) );
  SDFFRQX2TH out47_reg_0_ ( .D(n238), .SI(n1576), .SE(n1520), .CK(clk), .RN(
        n679), .Q(out47[0]) );
  SDFFRQX2TH out11_reg_0_ ( .D(n274), .SI(n2149), .SE(n1497), .CK(clk), .RN(
        n678), .Q(out11[0]) );
  SDFFRQX1TH out32_reg_1_ ( .D(n301), .SI(n1666), .SE(n1487), .CK(clk), .RN(
        n682), .Q(out32[1]) );
  SDFFRQX2TH out45_reg_0_ ( .D(n240), .SI(n2191), .SE(n1504), .CK(clk), .RN(
        n679), .Q(out45[0]) );
  SDFFRQX2TH out32_reg_0_ ( .D(n253), .SI(n2113), .SE(n1517), .CK(clk), .RN(
        n677), .Q(out32[0]) );
  SDFFRQX1TH out45_reg_4_ ( .D(n432), .SI(n1942), .SE(n1495), .CK(clk), .RN(
        n685), .Q(out45[4]) );
  SDFFRQX2TH count1_reg ( .D(n478), .SI(test_si), .SE(n1509), .CK(clk), .RN(
        n684), .Q(count1) );
  SDFFRQX1TH out47_reg_3_ ( .D(n382), .SI(n2262), .SE(n1496), .CK(clk), .RN(
        n683), .Q(out47[3]) );
  SDFFRQX2TH count2_reg_9_ ( .D(n498), .SI(count2[8]), .SE(n1505), .CK(clk), 
        .RN(n684), .Q(count2[9]) );
  SDFFRQX2TH count2_reg_1_ ( .D(n496), .SI(count2[0]), .SE(n1508), .CK(clk), 
        .RN(n684), .Q(count2[1]) );
  SDFFRQX2TH count2_reg_2_ ( .D(n495), .SI(count2[1]), .SE(n1468), .CK(clk), 
        .RN(n684), .Q(count2[2]) );
  SDFFRQX2TH count2_reg_3_ ( .D(n494), .SI(count2[2]), .SE(n1510), .CK(clk), 
        .RN(n683), .Q(count2[3]) );
  SDFFRQX2TH count2_reg_4_ ( .D(n493), .SI(count2[3]), .SE(n1510), .CK(clk), 
        .RN(n683), .Q(count2[4]) );
  SDFFRQX2TH count2_reg_5_ ( .D(n492), .SI(count2[4]), .SE(n1510), .CK(clk), 
        .RN(n683), .Q(count2[5]) );
  SDFFRQX2TH count2_reg_6_ ( .D(n491), .SI(count2[5]), .SE(n1505), .CK(clk), 
        .RN(n683), .Q(count2[6]) );
  SDFFRQX2TH count2_reg_7_ ( .D(n490), .SI(count2[6]), .SE(n1505), .CK(clk), 
        .RN(n683), .Q(count2[7]) );
  SDFFRQX2TH count2_reg_8_ ( .D(n489), .SI(count2[7]), .SE(n1505), .CK(clk), 
        .RN(n683), .Q(count2[8]) );
  SDFFRQX4TH count2_reg_0_ ( .D(n497), .SI(count1), .SE(n1508), .CK(clk), .RN(
        n685), .Q(count2[0]) );
  SDFFRXLTH out7_reg_4_ ( .D(n470), .SI(n2260), .SE(n1508), .CK(clk), .RN(
        reset), .Q(out7[4]), .QN(n1458) );
  SDFFRXLTH count_reg_7_ ( .D(n485), .SI(count[6]), .SE(n1508), .CK(clk), .RN(
        reset), .Q(count[7]), .QN(n1227) );
  SDFFRQX1TH out9_reg_3_ ( .D(n420), .SI(n1723), .SE(n1526), .CK(clk), .RN(
        n682), .Q(out9[3]) );
  SDFFRQX1TH out18_reg_3_ ( .D(n411), .SI(n1744), .SE(n1479), .CK(clk), .RN(
        n682), .Q(out18[3]) );
  SDFFRQX2TH out42_reg_1_ ( .D(n291), .SI(n2086), .SE(n1519), .CK(clk), .RN(
        n688), .Q(out42[1]) );
  SDFFRQX1TH out34_reg_3_ ( .D(n395), .SI(n1786), .SE(n1541), .CK(clk), .RN(
        n680), .Q(out34[3]) );
  AND4XLTH U3 ( .A(n1558), .B(n1555), .C(n1227), .D(n504), .Y(n594) );
  BUFX3TH U4 ( .A(n701), .Y(n675) );
  BUFX3TH U5 ( .A(n696), .Y(n684) );
  CLKBUFX1TH U8 ( .A(n594), .Y(n673) );
  CLKBUFX1TH U9 ( .A(n594), .Y(n672) );
  CLKBUFX1TH U10 ( .A(n672), .Y(n670) );
  CLKBUFX1TH U11 ( .A(n673), .Y(n669) );
  CLKBUFX1TH U12 ( .A(n673), .Y(n668) );
  CLKBUFX1TH U13 ( .A(n672), .Y(n671) );
  CLKBUFX1TH U14 ( .A(n671), .Y(n657) );
  CLKBUFX1TH U15 ( .A(n670), .Y(n658) );
  CLKBUFX1TH U16 ( .A(n668), .Y(n667) );
  CLKBUFX1TH U17 ( .A(n668), .Y(n666) );
  CLKBUFX1TH U18 ( .A(n670), .Y(n660) );
  CLKBUFX1TH U19 ( .A(n670), .Y(n659) );
  CLKBUFX1TH U20 ( .A(n672), .Y(n661) );
  CLKBUFX1TH U21 ( .A(n669), .Y(n662) );
  CLKBUFX1TH U22 ( .A(n669), .Y(n663) );
  CLKBUFX1TH U23 ( .A(n669), .Y(n664) );
  CLKBUFX1TH U24 ( .A(n681), .Y(n704) );
  CLKBUFX1TH U25 ( .A(n671), .Y(n656) );
  CLKBUFX1TH U26 ( .A(reset), .Y(n674) );
  CLKBUFX1TH U27 ( .A(n668), .Y(n665) );
  CLKBUFX1TH U28 ( .A(n674), .Y(n703) );
  CLKBUFX1TH U29 ( .A(n671), .Y(n655) );
  INVX2TH U30 ( .A(n597), .Y(n1225) );
  INVXLTH U31 ( .A(out10[0]), .Y(n1288) );
  INVXLTH U32 ( .A(out9[0]), .Y(n1287) );
  CLKBUFX1TH U33 ( .A(n665), .Y(n622) );
  INVXLTH U34 ( .A(out25[1]), .Y(n1388) );
  INVXLTH U35 ( .A(out5[1]), .Y(n1372) );
  INVXLTH U36 ( .A(out40[1]), .Y(n1402) );
  INVXLTH U37 ( .A(out37[1]), .Y(n1400) );
  INVXLTH U38 ( .A(out10[1]), .Y(n1376) );
  INVXLTH U39 ( .A(out9[1]), .Y(n1375) );
  INVXLTH U40 ( .A(out31[1]), .Y(n1394) );
  INVXLTH U41 ( .A(out44[1]), .Y(n1453) );
  INVXLTH U42 ( .A(out43[1]), .Y(n1405) );
  INVXLTH U43 ( .A(out6[4]), .Y(n1413) );
  INVXLTH U44 ( .A(out38[4]), .Y(n1443) );
  INVXLTH U45 ( .A(out5[4]), .Y(n1412) );
  INVXLTH U46 ( .A(out25[4]), .Y(n1430) );
  INVXLTH U47 ( .A(out2[4]), .Y(n1409) );
  INVXLTH U48 ( .A(out30[4]), .Y(n1435) );
  INVXLTH U49 ( .A(out33[4]), .Y(n1438) );
  INVXLTH U50 ( .A(out22[4]), .Y(n1427) );
  INVXLTH U51 ( .A(out26[4]), .Y(n1431) );
  INVXLTH U52 ( .A(out44[4]), .Y(n1449) );
  INVXLTH U53 ( .A(out21[4]), .Y(n1426) );
  INVXLTH U54 ( .A(out34[4]), .Y(n1439) );
  INVXLTH U55 ( .A(out15[4]), .Y(n1421) );
  INVXLTH U56 ( .A(out46[4]), .Y(n1451) );
  INVXLTH U57 ( .A(out9[4]), .Y(n1415) );
  INVXLTH U58 ( .A(out41[4]), .Y(n1446) );
  INVXLTH U59 ( .A(out40[4]), .Y(n1445) );
  CLKBUFX2TH U60 ( .A(n659), .Y(n642) );
  INVXLTH U61 ( .A(out43[4]), .Y(n1448) );
  INVXLTH U62 ( .A(out42[4]), .Y(n1447) );
  INVXLTH U63 ( .A(out24[4]), .Y(n1429) );
  INVXLTH U64 ( .A(out23[4]), .Y(n1428) );
  INVXLTH U65 ( .A(out37[4]), .Y(n1442) );
  INVXLTH U66 ( .A(out29[4]), .Y(n1434) );
  INVXLTH U67 ( .A(out17[4]), .Y(n1457) );
  INVXLTH U68 ( .A(out10[4]), .Y(n1416) );
  INVXLTH U69 ( .A(out0[3]), .Y(n1229) );
  INVXLTH U70 ( .A(out12[3]), .Y(n1241) );
  INVXLTH U71 ( .A(out33[3]), .Y(n1262) );
  INVXLTH U72 ( .A(out32[3]), .Y(n1261) );
  INVXLTH U73 ( .A(out16[3]), .Y(n1245) );
  INVXLTH U74 ( .A(out11[3]), .Y(n1240) );
  INVXLTH U75 ( .A(out10[3]), .Y(n1239) );
  INVXLTH U76 ( .A(out9[3]), .Y(n1238) );
  INVXLTH U77 ( .A(out8[3]), .Y(n1237) );
  INVXLTH U78 ( .A(out1[3]), .Y(n1230) );
  INVXLTH U79 ( .A(out46[3]), .Y(n1275) );
  INVXLTH U80 ( .A(out45[3]), .Y(n1274) );
  INVXLTH U81 ( .A(out44[3]), .Y(n1273) );
  INVXLTH U82 ( .A(out43[3]), .Y(n1272) );
  INVXLTH U83 ( .A(out42[3]), .Y(n1271) );
  INVXLTH U84 ( .A(out41[3]), .Y(n1270) );
  INVXLTH U85 ( .A(out40[3]), .Y(n1269) );
  INVXLTH U86 ( .A(out39[3]), .Y(n1268) );
  INVXLTH U87 ( .A(out38[3]), .Y(n1267) );
  INVXLTH U88 ( .A(out37[3]), .Y(n1266) );
  INVXLTH U89 ( .A(out34[3]), .Y(n1263) );
  INVXLTH U90 ( .A(out31[3]), .Y(n1260) );
  CLKBUFX2TH U91 ( .A(n657), .Y(n648) );
  INVXLTH U92 ( .A(out29[3]), .Y(n1258) );
  INVXLTH U93 ( .A(out30[3]), .Y(n1259) );
  INVXLTH U94 ( .A(out26[3]), .Y(n1255) );
  INVXLTH U95 ( .A(out25[3]), .Y(n1254) );
  INVXLTH U96 ( .A(out23[3]), .Y(n1252) );
  INVXLTH U97 ( .A(out24[3]), .Y(n1253) );
  INVXLTH U98 ( .A(out22[3]), .Y(n1251) );
  INVXLTH U99 ( .A(out21[3]), .Y(n1250) );
  INVXLTH U100 ( .A(out17[3]), .Y(n1246) );
  INVXLTH U101 ( .A(out15[3]), .Y(n1244) );
  CLKBUFX2TH U102 ( .A(n658), .Y(n644) );
  INVXLTH U103 ( .A(out7[3]), .Y(n1236) );
  INVXLTH U104 ( .A(out6[3]), .Y(n1235) );
  INVXLTH U105 ( .A(out5[3]), .Y(n1234) );
  INVXLTH U106 ( .A(out2[3]), .Y(n1231) );
  CLKBUFX2TH U107 ( .A(n656), .Y(n649) );
  INVXLTH U108 ( .A(out35[3]), .Y(n1264) );
  INVXLTH U109 ( .A(out36[3]), .Y(n1265) );
  INVX3TH U110 ( .A(n629), .Y(n602) );
  CLKBUFX2TH U111 ( .A(n657), .Y(n647) );
  INVXLTH U112 ( .A(out28[3]), .Y(n1257) );
  INVXLTH U113 ( .A(out27[3]), .Y(n1256) );
  INVXLTH U114 ( .A(out20[3]), .Y(n1249) );
  CLKBUFX2TH U115 ( .A(n657), .Y(n646) );
  INVXLTH U116 ( .A(out19[3]), .Y(n1248) );
  INVXLTH U117 ( .A(out18[3]), .Y(n1247) );
  INVX3TH U118 ( .A(n627), .Y(n604) );
  CLKBUFX2TH U119 ( .A(n658), .Y(n643) );
  INVXLTH U120 ( .A(out4[3]), .Y(n1233) );
  INVXLTH U121 ( .A(out3[3]), .Y(n1232) );
  CLKBUFX1TH U122 ( .A(n703), .Y(n697) );
  CLKBUFX2TH U123 ( .A(n658), .Y(n645) );
  INVXLTH U124 ( .A(out14[3]), .Y(n1243) );
  INVXLTH U125 ( .A(out13[3]), .Y(n1242) );
  CLKBUFX1TH U126 ( .A(n666), .Y(n619) );
  CLKBUFX1TH U127 ( .A(n666), .Y(n618) );
  CLKBUFX1TH U128 ( .A(n667), .Y(n616) );
  CLKBUFX1TH U129 ( .A(n667), .Y(n617) );
  INVXLTH U130 ( .A(out11[0]), .Y(n1289) );
  INVXLTH U131 ( .A(out34[0]), .Y(n1310) );
  INVXLTH U132 ( .A(out23[0]), .Y(n1299) );
  INVXLTH U133 ( .A(out41[0]), .Y(n1317) );
  CLKBUFX1TH U134 ( .A(n666), .Y(n620) );
  INVXLTH U135 ( .A(out37[0]), .Y(n1313) );
  INVX3TH U136 ( .A(n623), .Y(n608) );
  INVXLTH U137 ( .A(out2[0]), .Y(n1280) );
  INVXLTH U138 ( .A(out11[1]), .Y(n1459) );
  INVXLTH U139 ( .A(out26[1]), .Y(n1389) );
  INVXLTH U140 ( .A(out38[1]), .Y(n1452) );
  CLKBUFX2TH U141 ( .A(n661), .Y(n634) );
  INVXLTH U142 ( .A(out6[1]), .Y(n1373) );
  CLKBUFX2TH U143 ( .A(n664), .Y(n635) );
  INVXLTH U144 ( .A(out34[1]), .Y(n1397) );
  INVX3TH U145 ( .A(n621), .Y(n610) );
  INVXLTH U146 ( .A(out23[1]), .Y(n1386) );
  INVX3TH U147 ( .A(n618), .Y(n613) );
  INVXLTH U148 ( .A(out2[1]), .Y(n1369) );
  INVX3TH U149 ( .A(n619), .Y(n612) );
  INVX3TH U150 ( .A(n620), .Y(n611) );
  CLKBUFX2TH U151 ( .A(n669), .Y(n636) );
  INVXLTH U152 ( .A(out41[1]), .Y(n1403) );
  CLKBUFX2TH U153 ( .A(n660), .Y(n639) );
  CLKBUFX2TH U154 ( .A(n659), .Y(n641) );
  INVXLTH U155 ( .A(out35[4]), .Y(n1440) );
  INVXLTH U156 ( .A(out11[4]), .Y(n1417) );
  NAND2X3TH U157 ( .A(out0[4]), .B(n619), .Y(n597) );
  CLKBUFX2TH U158 ( .A(n660), .Y(n637) );
  INVX3TH U159 ( .A(n625), .Y(n606) );
  CLKBUFX2TH U160 ( .A(n660), .Y(n638) );
  INVXLTH U161 ( .A(out18[4]), .Y(n1423) );
  CLKBUFX1TH U162 ( .A(n701), .Y(n695) );
  INVX3TH U163 ( .A(n626), .Y(n605) );
  CLKBUFX2TH U164 ( .A(n659), .Y(n640) );
  INVXLTH U165 ( .A(out31[4]), .Y(n1436) );
  CLKBUFX1TH U166 ( .A(n692), .Y(n694) );
  INVX3TH U167 ( .A(n624), .Y(n607) );
  INVXLTH U168 ( .A(out3[4]), .Y(n1410) );
  CLKBUFX1TH U169 ( .A(n702), .Y(n700) );
  INVX3TH U170 ( .A(n622), .Y(n609) );
  INVXLTH U171 ( .A(out26[0]), .Y(n1302) );
  INVX3TH U172 ( .A(n628), .Y(n603) );
  CLKBUFX2TH U173 ( .A(n661), .Y(n633) );
  INVXLTH U174 ( .A(out44[2]), .Y(n1365) );
  INVXLTH U175 ( .A(out43[2]), .Y(n1364) );
  INVXLTH U176 ( .A(out42[2]), .Y(n1363) );
  CLKBUFX1TH U177 ( .A(n662), .Y(n632) );
  INVXLTH U178 ( .A(out41[2]), .Y(n1362) );
  INVXLTH U179 ( .A(out40[2]), .Y(n1361) );
  CLKBUFX1TH U180 ( .A(n662), .Y(n631) );
  INVXLTH U181 ( .A(out39[2]), .Y(n1360) );
  INVXLTH U182 ( .A(out38[2]), .Y(n1359) );
  CLKBUFX1TH U183 ( .A(n662), .Y(n630) );
  INVXLTH U184 ( .A(out37[2]), .Y(n1358) );
  INVXLTH U185 ( .A(out36[2]), .Y(n1357) );
  CLKBUFX1TH U186 ( .A(n663), .Y(n629) );
  INVX3TH U187 ( .A(n617), .Y(n614) );
  INVXLTH U188 ( .A(out35[2]), .Y(n1356) );
  INVXLTH U189 ( .A(out34[2]), .Y(n1355) );
  CLKBUFX1TH U190 ( .A(n663), .Y(n628) );
  INVXLTH U191 ( .A(out33[2]), .Y(n1354) );
  CLKBUFX1TH U192 ( .A(n663), .Y(n627) );
  INVXLTH U193 ( .A(out31[2]), .Y(n1352) );
  INVXLTH U194 ( .A(out30[2]), .Y(n1351) );
  CLKBUFX1TH U195 ( .A(n664), .Y(n626) );
  INVXLTH U196 ( .A(out29[2]), .Y(n1350) );
  CLKBUFX1TH U197 ( .A(n664), .Y(n625) );
  INVXLTH U198 ( .A(out27[2]), .Y(n1348) );
  INVXLTH U199 ( .A(out26[2]), .Y(n1460) );
  CLKBUFX1TH U200 ( .A(n664), .Y(n624) );
  INVXLTH U201 ( .A(out25[2]), .Y(n1347) );
  CLKBUFX1TH U202 ( .A(n704), .Y(n693) );
  INVXLTH U203 ( .A(out24[2]), .Y(n1346) );
  CLKBUFX1TH U204 ( .A(n665), .Y(n623) );
  INVXLTH U205 ( .A(out23[2]), .Y(n1345) );
  INVXLTH U206 ( .A(out22[2]), .Y(n1344) );
  INVXLTH U207 ( .A(out21[2]), .Y(n1343) );
  INVXLTH U208 ( .A(out20[2]), .Y(n1342) );
  INVXLTH U209 ( .A(out19[2]), .Y(n1341) );
  INVXLTH U210 ( .A(out18[2]), .Y(n1340) );
  INVX3TH U211 ( .A(n632), .Y(n599) );
  INVXLTH U212 ( .A(out17[2]), .Y(n1339) );
  INVXLTH U213 ( .A(out16[2]), .Y(n1338) );
  INVXLTH U214 ( .A(out15[2]), .Y(n1337) );
  CLKBUFX2TH U215 ( .A(n655), .Y(n653) );
  INVXLTH U216 ( .A(out13[2]), .Y(n1335) );
  INVXLTH U217 ( .A(out11[2]), .Y(n1333) );
  CLKBUFX1TH U218 ( .A(n704), .Y(n692) );
  INVXLTH U219 ( .A(out10[2]), .Y(n1332) );
  CLKBUFX1TH U220 ( .A(n703), .Y(n698) );
  INVXLTH U221 ( .A(out9[2]), .Y(n1331) );
  INVXLTH U222 ( .A(out8[2]), .Y(n1330) );
  CLKBUFX2TH U223 ( .A(n655), .Y(n652) );
  INVXLTH U224 ( .A(out7[2]), .Y(n1329) );
  INVXLTH U225 ( .A(out6[2]), .Y(n1328) );
  INVXLTH U226 ( .A(out5[2]), .Y(n1327) );
  INVXLTH U227 ( .A(out4[2]), .Y(n1326) );
  INVX3TH U228 ( .A(n631), .Y(n600) );
  INVXLTH U229 ( .A(out3[2]), .Y(n1325) );
  CLKBUFX2TH U230 ( .A(n656), .Y(n650) );
  INVXLTH U231 ( .A(out2[2]), .Y(n1324) );
  INVX3TH U232 ( .A(n630), .Y(n601) );
  CLKBUFX2TH U233 ( .A(n656), .Y(n651) );
  INVXLTH U234 ( .A(out1[2]), .Y(n1323) );
  CLKBUFX1TH U235 ( .A(n674), .Y(n702) );
  CLKBUFX1TH U236 ( .A(n665), .Y(n621) );
  INVXLTH U237 ( .A(out0[2]), .Y(n1321) );
  CLKBUFX1TH U238 ( .A(n702), .Y(n699) );
  INVX3TH U239 ( .A(n661), .Y(n598) );
  INVX3TH U240 ( .A(n616), .Y(n615) );
  INVXLTH U241 ( .A(out46[2]), .Y(n1367) );
  INVXLTH U242 ( .A(count[8]), .Y(n1228) );
  CLKBUFX1TH U243 ( .A(n703), .Y(n696) );
  INVXLTH U244 ( .A(count[9]), .Y(n1226) );
  CLKBUFX2TH U245 ( .A(n655), .Y(n654) );
  OAI22XLTH U246 ( .A0(n607), .A1(n2219), .B0(n668), .B1(n1978), .Y(n470) );
  AO22XLTH U247 ( .A0(count2[8]), .A1(n597), .B0(N23), .B1(n1225), .Y(n489) );
  AO22XLTH U248 ( .A0(count2[7]), .A1(n597), .B0(N22), .B1(n1225), .Y(n490) );
  AO22XLTH U249 ( .A0(count2[6]), .A1(n597), .B0(N21), .B1(n1225), .Y(n491) );
  AO22XLTH U250 ( .A0(count2[5]), .A1(n597), .B0(N20), .B1(n1225), .Y(n492) );
  AO22XLTH U251 ( .A0(count2[4]), .A1(n597), .B0(N19), .B1(n1225), .Y(n493) );
  AO22XLTH U252 ( .A0(count2[3]), .A1(n597), .B0(N18), .B1(n1225), .Y(n494) );
  AO22XLTH U253 ( .A0(count2[2]), .A1(n597), .B0(N17), .B1(n1225), .Y(n495) );
  AO22XLTH U254 ( .A0(count2[1]), .A1(n597), .B0(N16), .B1(n1225), .Y(n496) );
  AO22XLTH U255 ( .A0(count2[9]), .A1(n597), .B0(N24), .B1(n1225), .Y(n498) );
  OAI2BB2XLTH U256 ( .B0(n598), .B1(n1571), .A0N(out47[3]), .A1N(n615), .Y(
        n382) );
  OAI22XLTH U257 ( .A0(n604), .A1(n2192), .B0(n642), .B1(n2098), .Y(n432) );
  OAI22XLTH U258 ( .A0(n608), .A1(n1664), .B0(n646), .B1(n1666), .Y(n253) );
  OAI22XLTH U259 ( .A0(n607), .A1(n1592), .B0(n622), .B1(n1594), .Y(n240) );
  OAI22XLTH U260 ( .A0(n611), .A1(n2228), .B0(n624), .B1(n2068), .Y(n301) );
  OAI22XLTH U261 ( .A0(n610), .A1(n1976), .B0(n670), .B1(n1837), .Y(n274) );
  OAI2BB2XLTH U262 ( .B0(n598), .B1(n1565), .A0N(out47[0]), .A1N(n615), .Y(
        n238) );
  OAI22XLTH U263 ( .A0(n608), .A1(n1685), .B0(n661), .B1(n1828), .Y(n244) );
  OAI22XLTH U264 ( .A0(n609), .A1(n1625), .B0(n643), .B1(n1696), .Y(n269) );
  OAI22XLTH U265 ( .A0(n611), .A1(n1643), .B0(n622), .B1(n1831), .Y(n262) );
  OAI22XLTH U266 ( .A0(n610), .A1(n1613), .B0(n657), .B1(n1972), .Y(n276) );
  OAI22XLTH U267 ( .A0(n608), .A1(n1676), .B0(n673), .B1(n1825), .Y(n248) );
  OAI22XLTH U268 ( .A0(n608), .A1(n1670), .B0(n638), .B1(n1834), .Y(n251) );
  OAI22XLTH U269 ( .A0(n610), .A1(n1973), .B0(n643), .B1(n1975), .Y(n275) );
  OAI22XLTH U270 ( .A0(n610), .A1(n1598), .B0(n635), .B1(n1822), .Y(n283) );
  OAI22XLTH U271 ( .A0(n613), .A1(n2234), .B0(n650), .B1(n2146), .Y(n322) );
  OAI2BB2XLTH U272 ( .B0(n598), .B1(n1574), .A0N(n1553), .A1N(n615), .Y(n286)
         );
  OAI2B2XLTH U273 ( .A1N(in[1]), .A0(n598), .B0(n2257), .B1(n622), .Y(n333) );
  OAI22XLTH U274 ( .A0(n610), .A1(n2225), .B0(n636), .B1(n2107), .Y(n288) );
  OAI22XLTH U275 ( .A0(n612), .A1(n2048), .B0(n660), .B1(n2104), .Y(n312) );
  OAI22XLTH U276 ( .A0(n613), .A1(n2036), .B0(n651), .B1(n2101), .Y(n317) );
  OAI22XLTH U277 ( .A0(n612), .A1(n2246), .B0(n655), .B1(n2143), .Y(n307) );
  OAI22XLTH U278 ( .A0(n612), .A1(n2054), .B0(n616), .B1(n2245), .Y(n308) );
  OAI22XLTH U279 ( .A0(n611), .A1(n2237), .B0(n635), .B1(n2140), .Y(n295) );
  OAI22XLTH U280 ( .A0(n613), .A1(n2243), .B0(n634), .B1(n2137), .Y(n327) );
  OAI22XLTH U281 ( .A0(n613), .A1(n2018), .B0(n634), .B1(n2242), .Y(n328) );
  OAI22XLTH U282 ( .A0(n611), .A1(n2081), .B0(n636), .B1(n2239), .Y(n293) );
  OAI22XLTH U283 ( .A0(n611), .A1(n2084), .B0(n636), .B1(n2221), .Y(n290) );
  OAI22XLTH U284 ( .A0(n611), .A1(n2240), .B0(n636), .B1(n2125), .Y(n292) );
  OAI22XLTH U285 ( .A0(n611), .A1(n2078), .B0(n635), .B1(n2236), .Y(n296) );
  OAI22XLTH U286 ( .A0(n611), .A1(n2072), .B0(n635), .B1(n2134), .Y(n299) );
  OAI22XLTH U287 ( .A0(n612), .A1(n2051), .B0(n667), .B1(n2131), .Y(n310) );
  OAI22XLTH U288 ( .A0(n613), .A1(n2231), .B0(n634), .B1(n2233), .Y(n323) );
  OAI22XLTH U289 ( .A0(n613), .A1(n2024), .B0(n634), .B1(n2230), .Y(n324) );
  OAI22XLTH U290 ( .A0(n614), .A1(n2012), .B0(n633), .B1(n2128), .Y(n331) );
  OAI22XLTH U291 ( .A0(n612), .A1(n2066), .B0(n667), .B1(n2227), .Y(n302) );
  OAI22XLTH U292 ( .A0(n611), .A1(n2222), .B0(n636), .B1(n2224), .Y(n289) );
  OAI2BB2XLTH U293 ( .B0(n598), .B1(n1577), .A0N(out47[4]), .A1N(n615), .Y(
        n430) );
  OAI22XLTH U294 ( .A0(n605), .A1(n2204), .B0(n640), .B1(n2113), .Y(n446) );
  OAI22XLTH U295 ( .A0(n606), .A1(n2183), .B0(n638), .B1(n2089), .Y(n461) );
  OAI22XLTH U296 ( .A0(n605), .A1(n2159), .B0(n641), .B1(n2215), .Y(n439) );
  OAI22XLTH U297 ( .A0(n599), .A1(n2207), .B0(n634), .B1(n2110), .Y(n474) );
  OAI22XLTH U298 ( .A0(n607), .A1(n2213), .B0(n629), .B1(n2218), .Y(n471) );
  OAI22XLTH U299 ( .A0(n605), .A1(n2210), .B0(n644), .B1(n2194), .Y(n451) );
  OAI22XLTH U300 ( .A0(n605), .A1(n2201), .B0(n640), .B1(n2185), .Y(n443) );
  OAI22XLTH U301 ( .A0(n605), .A1(n2216), .B0(n641), .B1(n2095), .Y(n438) );
  OAI22XLTH U302 ( .A0(n607), .A1(n1982), .B0(n627), .B1(n2212), .Y(n472) );
  OAI22XLTH U303 ( .A0(n606), .A1(n2165), .B0(n639), .B1(n2209), .Y(n452) );
  OAI22XLTH U304 ( .A0(n607), .A1(n1561), .B0(n633), .B1(n2206), .Y(n475) );
  OAI22XLTH U305 ( .A0(n607), .A1(n2180), .B0(n637), .B1(n2149), .Y(n467) );
  OAI22XLTH U306 ( .A0(n606), .A1(n2198), .B0(n639), .B1(n2161), .Y(n454) );
  OAI22XLTH U307 ( .A0(n605), .A1(n2156), .B0(n640), .B1(n2203), .Y(n447) );
  OAI22XLTH U308 ( .A0(n605), .A1(n2006), .B0(n640), .B1(n2200), .Y(n444) );
  OAI22XLTH U309 ( .A0(n606), .A1(n2090), .B0(n638), .B1(n2152), .Y(n460) );
  OAI22XLTH U310 ( .A0(n606), .A1(n2189), .B0(n639), .B1(n2197), .Y(n455) );
  OAI22XLTH U311 ( .A0(n605), .A1(n2195), .B0(n639), .B1(n2092), .Y(n450) );
  OAI22XLTH U312 ( .A0(n604), .A1(n2171), .B0(n642), .B1(n2191), .Y(n433) );
  OAI22XLTH U313 ( .A0(n606), .A1(n2000), .B0(n638), .B1(n2188), .Y(n456) );
  OAI22XLTH U314 ( .A0(n605), .A1(n2186), .B0(n641), .B1(n2122), .Y(n442) );
  OAI22XLTH U315 ( .A0(n606), .A1(n1994), .B0(n637), .B1(n2182), .Y(n462) );
  OAI22XLTH U316 ( .A0(n604), .A1(n2099), .B0(n642), .B1(n1576), .Y(n431) );
  OAI22XLTH U317 ( .A0(n607), .A1(n1985), .B0(n626), .B1(n2179), .Y(n468) );
  OAI22XLTH U318 ( .A0(n604), .A1(n2177), .B0(n642), .B1(n2167), .Y(n435) );
  OAI22XLTH U319 ( .A0(n604), .A1(n2096), .B0(n641), .B1(n2173), .Y(n437) );
  OAI22XLTH U320 ( .A0(n604), .A1(n2174), .B0(n642), .B1(n2176), .Y(n436) );
  OAI22XLTH U321 ( .A0(n604), .A1(n2168), .B0(n642), .B1(n2170), .Y(n434) );
  OAI22XLTH U322 ( .A0(n606), .A1(n2162), .B0(n639), .B1(n2164), .Y(n453) );
  OAI22XLTH U323 ( .A0(n605), .A1(n2009), .B0(n641), .B1(n2158), .Y(n440) );
  OAI22XLTH U324 ( .A0(n605), .A1(n2003), .B0(n640), .B1(n2155), .Y(n448) );
  OAI22XLTH U325 ( .A0(n606), .A1(n2153), .B0(n638), .B1(n2116), .Y(n459) );
  OAI22XLTH U326 ( .A0(n607), .A1(n2150), .B0(n637), .B1(n2119), .Y(n466) );
  OAI22XLTH U327 ( .A0(n601), .A1(n1940), .B0(n650), .B1(n1942), .Y(n384) );
  OAI22XLTH U328 ( .A0(n603), .A1(n1883), .B0(n645), .B1(n1960), .Y(n413) );
  OAI22XLTH U329 ( .A0(n603), .A1(n1958), .B0(n645), .B1(n1969), .Y(n417) );
  OAI2B2XLTH U330 ( .A1N(in[3]), .A0(n598), .B0(n2254), .B1(n621), .Y(n429) );
  OAI22XLTH U331 ( .A0(n602), .A1(n1904), .B0(n647), .B1(n1861), .Y(n402) );
  OAI22XLTH U332 ( .A0(n604), .A1(n2255), .B0(n643), .B1(n1945), .Y(n428) );
  OAI22XLTH U333 ( .A0(n602), .A1(n1913), .B0(n648), .B1(n1963), .Y(n397) );
  OAI22XLTH U334 ( .A0(n603), .A1(n1970), .B0(n645), .B1(n1840), .Y(n416) );
  OAI22XLTH U335 ( .A0(n603), .A1(n2261), .B0(n644), .B1(n1948), .Y(n421) );
  OAI22XLTH U336 ( .A0(n615), .A1(n1781), .B0(n627), .B1(n1690), .Y(n349) );
  OAI22XLTH U337 ( .A0(n614), .A1(n1817), .B0(n633), .B1(n1693), .Y(n336) );
  OAI22XLTH U338 ( .A0(n601), .A1(n1928), .B0(n649), .B1(n1930), .Y(n388) );
  OAI22XLTH U339 ( .A0(n601), .A1(n1868), .B0(n649), .B1(n1918), .Y(n392) );
  OAI22XLTH U340 ( .A0(n602), .A1(n1967), .B0(n648), .B1(n1915), .Y(n395) );
  OAI22XLTH U341 ( .A0(n602), .A1(n1964), .B0(n648), .B1(n1966), .Y(n396) );
  OAI22XLTH U342 ( .A0(n602), .A1(n1865), .B0(n647), .B1(n1909), .Y(n400) );
  OAI22XLTH U343 ( .A0(n602), .A1(n1892), .B0(n646), .B1(n1897), .Y(n406) );
  OAI22XLTH U344 ( .A0(n603), .A1(n1961), .B0(n645), .B1(n1885), .Y(n412) );
  OAI22XLTH U345 ( .A0(n603), .A1(n1955), .B0(n644), .B1(n1957), .Y(n418) );
  OAI22XLTH U346 ( .A0(n603), .A1(n1952), .B0(n644), .B1(n1954), .Y(n419) );
  OAI22XLTH U347 ( .A0(n603), .A1(n1949), .B0(n644), .B1(n1951), .Y(n420) );
  OAI22XLTH U348 ( .A0(n604), .A1(n1946), .B0(n643), .B1(n1873), .Y(n427) );
  OAI22XLTH U349 ( .A0(n601), .A1(n1943), .B0(n650), .B1(n1570), .Y(n383) );
  OAI22XLTH U350 ( .A0(n601), .A1(n1937), .B0(n650), .B1(n1939), .Y(n385) );
  OAI22XLTH U351 ( .A0(n601), .A1(n1934), .B0(n650), .B1(n1936), .Y(n386) );
  OAI22XLTH U352 ( .A0(n601), .A1(n1931), .B0(n650), .B1(n1933), .Y(n387) );
  OAI22XLTH U353 ( .A0(n601), .A1(n1925), .B0(n649), .B1(n1927), .Y(n389) );
  OAI22XLTH U354 ( .A0(n601), .A1(n1922), .B0(n649), .B1(n1924), .Y(n390) );
  OAI22XLTH U355 ( .A0(n601), .A1(n1919), .B0(n649), .B1(n1921), .Y(n391) );
  OAI22XLTH U356 ( .A0(n601), .A1(n1916), .B0(n648), .B1(n1870), .Y(n394) );
  OAI22XLTH U357 ( .A0(n602), .A1(n1907), .B0(n648), .B1(n1912), .Y(n398) );
  OAI22XLTH U358 ( .A0(n602), .A1(n1910), .B0(n648), .B1(n1906), .Y(n399) );
  OAI22XLTH U359 ( .A0(n602), .A1(n1901), .B0(n647), .B1(n1903), .Y(n403) );
  OAI22XLTH U360 ( .A0(n602), .A1(n1895), .B0(n647), .B1(n1900), .Y(n404) );
  OAI22XLTH U361 ( .A0(n602), .A1(n1898), .B0(n647), .B1(n1894), .Y(n405) );
  OAI22XLTH U362 ( .A0(n602), .A1(n1889), .B0(n646), .B1(n1891), .Y(n407) );
  OAI22XLTH U363 ( .A0(n602), .A1(n1859), .B0(n646), .B1(n1888), .Y(n408) );
  OAI22XLTH U364 ( .A0(n603), .A1(n1886), .B0(n646), .B1(n1852), .Y(n411) );
  OAI22XLTH U365 ( .A0(n603), .A1(n1844), .B0(n645), .B1(n1882), .Y(n414) );
  OAI22XLTH U366 ( .A0(n604), .A1(n1880), .B0(n644), .B1(n2260), .Y(n422) );
  OAI22XLTH U367 ( .A0(n604), .A1(n1877), .B0(n643), .B1(n1879), .Y(n423) );
  OAI22XLTH U368 ( .A0(n604), .A1(n1850), .B0(n643), .B1(n1876), .Y(n424) );
  OAI22XLTH U369 ( .A0(n604), .A1(n1874), .B0(n643), .B1(n1846), .Y(n426) );
  OAI22XLTH U370 ( .A0(n601), .A1(n1871), .B0(n649), .B1(n1867), .Y(n393) );
  OAI22XLTH U371 ( .A0(n602), .A1(n1862), .B0(n647), .B1(n1864), .Y(n401) );
  OAI22XLTH U372 ( .A0(n603), .A1(n1856), .B0(n646), .B1(n1858), .Y(n409) );
  CLKBUFX4TH U373 ( .A(n698), .Y(n681) );
  OAI22XLTH U374 ( .A0(n603), .A1(n1853), .B0(n646), .B1(n1855), .Y(n410) );
  CLKBUFX4TH U375 ( .A(n697), .Y(n683) );
  OAI22XLTH U376 ( .A0(n604), .A1(n1847), .B0(n643), .B1(n1849), .Y(n425) );
  CLKBUFX4TH U377 ( .A(n697), .Y(n682) );
  OAI22XLTH U378 ( .A0(n603), .A1(n1841), .B0(n645), .B1(n1843), .Y(n415) );
  OAI22XLTH U379 ( .A0(n608), .A1(n1673), .B0(n650), .B1(n1675), .Y(n249) );
  OAI22XLTH U380 ( .A0(n609), .A1(n1619), .B0(n637), .B1(n1621), .Y(n271) );
  OAI22XLTH U381 ( .A0(n609), .A1(n1616), .B0(n623), .B1(n1618), .Y(n272) );
  OAI22XLTH U382 ( .A0(n610), .A1(n2249), .B0(n637), .B1(n1597), .Y(n284) );
  OAI22XLTH U383 ( .A0(n613), .A1(n2030), .B0(n653), .B1(n2032), .Y(n319) );
  OAI22XLTH U384 ( .A0(n608), .A1(n1652), .B0(n638), .B1(n1654), .Y(n257) );
  OAI22XLTH U385 ( .A0(n609), .A1(n1634), .B0(n618), .B1(n1636), .Y(n265) );
  OAI22XLTH U386 ( .A0(n610), .A1(n1838), .B0(n654), .B1(n1615), .Y(n273) );
  OAI22XLTH U387 ( .A0(n610), .A1(n1589), .B0(n644), .B1(n1600), .Y(n281) );
  OAI22XLTH U388 ( .A0(n609), .A1(n1631), .B0(n621), .B1(n1633), .Y(n266) );
  OAI22XLTH U389 ( .A0(n609), .A1(n1820), .B0(n642), .B1(n1651), .Y(n258) );
  OAI22XLTH U390 ( .A0(n608), .A1(n1667), .B0(n642), .B1(n1669), .Y(n252) );
  OAI22XLTH U391 ( .A0(n610), .A1(n1610), .B0(n636), .B1(n1612), .Y(n277) );
  OAI22XLTH U392 ( .A0(n608), .A1(n1679), .B0(n651), .B1(n1681), .Y(n246) );
  OAI22XLTH U393 ( .A0(n608), .A1(n1835), .B0(n641), .B1(n1672), .Y(n250) );
  OAI22XLTH U394 ( .A0(n610), .A1(n1607), .B0(n649), .B1(n1609), .Y(n278) );
  OAI22XLTH U395 ( .A0(n609), .A1(n1628), .B0(n645), .B1(n1630), .Y(n267) );
  OAI22XLTH U396 ( .A0(n607), .A1(n1595), .B0(n631), .B1(n1564), .Y(n239) );
  OAI22XLTH U397 ( .A0(n608), .A1(n1655), .B0(n641), .B1(n1657), .Y(n256) );
  OAI22XLTH U398 ( .A0(n609), .A1(n1697), .B0(n633), .B1(n1627), .Y(n268) );
  OAI22XLTH U399 ( .A0(n609), .A1(n1832), .B0(n640), .B1(n1645), .Y(n261) );
  OAI22XLTH U400 ( .A0(n609), .A1(n1622), .B0(n634), .B1(n1624), .Y(n270) );
  OAI22XLTH U401 ( .A0(n609), .A1(n1640), .B0(n648), .B1(n1642), .Y(n263) );
  OAI22XLTH U402 ( .A0(n608), .A1(n1658), .B0(n640), .B1(n1660), .Y(n255) );
  OAI22XLTH U403 ( .A0(n607), .A1(n1829), .B0(n673), .B1(n2086), .Y(n243) );
  OAI22XLTH U404 ( .A0(n607), .A1(n2087), .B0(n639), .B1(n1687), .Y(n242) );
  OAI22XLTH U405 ( .A0(n610), .A1(n1601), .B0(n658), .B1(n1603), .Y(n280) );
  OAI22XLTH U406 ( .A0(n608), .A1(n1682), .B0(n653), .B1(n1684), .Y(n245) );
  OAI2B2XLTH U407 ( .A1N(in[0]), .A0(n598), .B0(n2248), .B1(n620), .Y(n285) );
  OAI22XLTH U408 ( .A0(n609), .A1(n1646), .B0(n620), .B1(n1648), .Y(n260) );
  OAI22XLTH U409 ( .A0(n608), .A1(n1826), .B0(n652), .B1(n1678), .Y(n247) );
  OAI22XLTH U410 ( .A0(n608), .A1(n1661), .B0(n644), .B1(n1663), .Y(n254) );
  CLKBUFX4TH U411 ( .A(n700), .Y(n676) );
  OAI22XLTH U412 ( .A0(n607), .A1(n1688), .B0(n654), .B1(n1591), .Y(n241) );
  CLKBUFX4TH U413 ( .A(n699), .Y(n678) );
  OAI22XLTH U414 ( .A0(n610), .A1(n1604), .B0(n672), .B1(n1606), .Y(n279) );
  OAI22XLTH U415 ( .A0(n609), .A1(n1637), .B0(n647), .B1(n1639), .Y(n264) );
  OAI22XLTH U416 ( .A0(n610), .A1(n1823), .B0(n632), .B1(n1588), .Y(n282) );
  OAI22XLTH U417 ( .A0(n612), .A1(n2057), .B0(n671), .B1(n2059), .Y(n305) );
  OAI22XLTH U418 ( .A0(n611), .A1(n2075), .B0(n635), .B1(n2077), .Y(n297) );
  OAI22XLTH U419 ( .A0(n614), .A1(n2258), .B0(n633), .B1(n2011), .Y(n332) );
  OAI22XLTH U420 ( .A0(n612), .A1(n2045), .B0(n659), .B1(n2047), .Y(n313) );
  OAI22XLTH U421 ( .A0(n613), .A1(n2147), .B0(n652), .B1(n2026), .Y(n321) );
  OAI22XLTH U422 ( .A0(n613), .A1(n2027), .B0(n649), .B1(n2029), .Y(n320) );
  OAI22XLTH U423 ( .A0(n612), .A1(n2042), .B0(n648), .B1(n2044), .Y(n314) );
  OAI22XLTH U424 ( .A0(n614), .A1(n2015), .B0(n633), .B1(n2017), .Y(n329) );
  OAI22XLTH U425 ( .A0(n612), .A1(n2144), .B0(n636), .B1(n2056), .Y(n306) );
  OAI22XLTH U426 ( .A0(n613), .A1(n2021), .B0(n634), .B1(n2023), .Y(n325) );
  OAI22XLTH U427 ( .A0(n611), .A1(n2141), .B0(n635), .B1(n2080), .Y(n294) );
  OAI22XLTH U428 ( .A0(n611), .A1(n2069), .B0(n665), .B1(n2071), .Y(n300) );
  OAI22XLTH U429 ( .A0(n613), .A1(n2138), .B0(n634), .B1(n2020), .Y(n326) );
  OAI22XLTH U430 ( .A0(n611), .A1(n2135), .B0(n635), .B1(n2074), .Y(n298) );
  OAI22XLTH U431 ( .A0(n612), .A1(n2039), .B0(n647), .B1(n2041), .Y(n315) );
  OAI22XLTH U432 ( .A0(n610), .A1(n2108), .B0(n656), .B1(n1573), .Y(n287) );
  OAI22XLTH U433 ( .A0(n612), .A1(n2060), .B0(n628), .B1(n2062), .Y(n304) );
  OAI22XLTH U434 ( .A0(n613), .A1(n2102), .B0(n646), .B1(n2038), .Y(n316) );
  OAI22XLTH U435 ( .A0(n612), .A1(n2132), .B0(n635), .B1(n2053), .Y(n309) );
  OAI22XLTH U436 ( .A0(n612), .A1(n2105), .B0(n645), .B1(n2050), .Y(n311) );
  OAI22XLTH U437 ( .A0(n613), .A1(n2033), .B0(n639), .B1(n2035), .Y(n318) );
  OAI22XLTH U438 ( .A0(n613), .A1(n2129), .B0(n633), .B1(n2014), .Y(n330) );
  OAI22XLTH U439 ( .A0(n612), .A1(n2063), .B0(n662), .B1(n2065), .Y(n303) );
  OAI22XLTH U440 ( .A0(n611), .A1(n2126), .B0(n636), .B1(n2083), .Y(n291) );
  OAI22XLTH U441 ( .A0(n606), .A1(n1991), .B0(n637), .B1(n1993), .Y(n463) );
  OAI22XLTH U442 ( .A0(n605), .A1(n2093), .B0(n639), .B1(n2002), .Y(n449) );
  OAI22XLTH U443 ( .A0(n605), .A1(n2123), .B0(n641), .B1(n2008), .Y(n441) );
  OAI22XLTH U444 ( .A0(n606), .A1(n2120), .B0(n637), .B1(n1987), .Y(n465) );
  OAI22XLTH U445 ( .A0(n606), .A1(n1997), .B0(n638), .B1(n1999), .Y(n457) );
  CLKBUFX4TH U446 ( .A(n694), .Y(n688) );
  OAI22XLTH U447 ( .A0(n606), .A1(n1988), .B0(n637), .B1(n1990), .Y(n464) );
  CLKBUFX4TH U448 ( .A(n695), .Y(n687) );
  OAI22XLTH U449 ( .A0(n606), .A1(n2117), .B0(n638), .B1(n1996), .Y(n458) );
  CLKBUFX4TH U450 ( .A(n695), .Y(n686) );
  OAI22XLTH U451 ( .A0(n605), .A1(n2114), .B0(n640), .B1(n2005), .Y(n445) );
  OAI22XLTH U452 ( .A0(n607), .A1(n1979), .B0(n625), .B1(n1984), .Y(n469) );
  OAI22XLTH U453 ( .A0(n607), .A1(n2111), .B0(n663), .B1(n1981), .Y(n473) );
  OAI22XLTH U454 ( .A0(n615), .A1(n1772), .B0(n625), .B1(n1585), .Y(n353) );
  OAI22XLTH U455 ( .A0(n600), .A1(n1733), .B0(n652), .B1(n1582), .Y(n367) );
  OAI22XLTH U456 ( .A0(n600), .A1(n1730), .B0(n652), .B1(n1579), .Y(n369) );
  CLKBUFX4TH U457 ( .A(n700), .Y(n677) );
  OAI22XLTH U458 ( .A0(n609), .A1(n1649), .B0(n617), .B1(n1819), .Y(n259) );
  OAI22XLTH U459 ( .A0(n603), .A1(n1766), .B0(n624), .B1(n1768), .Y(n355) );
  OAI22XLTH U460 ( .A0(n614), .A1(n1694), .B0(n633), .B1(n1567), .Y(n335) );
  OAI22XLTH U461 ( .A0(n614), .A1(n1814), .B0(n666), .B1(n1816), .Y(n337) );
  OAI22XLTH U462 ( .A0(n614), .A1(n1811), .B0(n619), .B1(n1813), .Y(n338) );
  OAI22XLTH U463 ( .A0(n614), .A1(n1808), .B0(n632), .B1(n1810), .Y(n339) );
  OAI22XLTH U464 ( .A0(n614), .A1(n1805), .B0(n632), .B1(n1807), .Y(n340) );
  OAI22XLTH U465 ( .A0(n614), .A1(n1802), .B0(n631), .B1(n1804), .Y(n341) );
  OAI22XLTH U466 ( .A0(n614), .A1(n1799), .B0(n631), .B1(n1801), .Y(n342) );
  CLKBUFX4TH U467 ( .A(n693), .Y(n689) );
  OAI22XLTH U468 ( .A0(n614), .A1(n1796), .B0(n630), .B1(n1798), .Y(n343) );
  OAI22XLTH U469 ( .A0(n614), .A1(n1793), .B0(n630), .B1(n1795), .Y(n344) );
  OAI22XLTH U470 ( .A0(n615), .A1(n1790), .B0(n629), .B1(n1792), .Y(n345) );
  OAI22XLTH U471 ( .A0(n614), .A1(n1787), .B0(n629), .B1(n1789), .Y(n346) );
  OAI22XLTH U472 ( .A0(n615), .A1(n1784), .B0(n628), .B1(n1786), .Y(n347) );
  OAI22XLTH U473 ( .A0(n615), .A1(n1691), .B0(n628), .B1(n1783), .Y(n348) );
  OAI22XLTH U474 ( .A0(n615), .A1(n1778), .B0(n627), .B1(n1780), .Y(n350) );
  OAI22XLTH U475 ( .A0(n615), .A1(n1775), .B0(n626), .B1(n1777), .Y(n351) );
  OAI22XLTH U476 ( .A0(n615), .A1(n1586), .B0(n626), .B1(n1774), .Y(n352) );
  OAI22XLTH U477 ( .A0(n615), .A1(n1769), .B0(n625), .B1(n1771), .Y(n354) );
  OAI22XLTH U478 ( .A0(n599), .A1(n1763), .B0(n624), .B1(n1765), .Y(n356) );
  CLKBUFX4TH U479 ( .A(n693), .Y(n690) );
  OAI22XLTH U480 ( .A0(n599), .A1(n1760), .B0(n623), .B1(n1762), .Y(n357) );
  OAI22XLTH U481 ( .A0(n599), .A1(n1757), .B0(n623), .B1(n1759), .Y(n358) );
  OAI22XLTH U482 ( .A0(n599), .A1(n1754), .B0(n630), .B1(n1756), .Y(n359) );
  OAI22XLTH U483 ( .A0(n599), .A1(n1751), .B0(n654), .B1(n1753), .Y(n360) );
  OAI22XLTH U484 ( .A0(n599), .A1(n1748), .B0(n653), .B1(n1750), .Y(n361) );
  OAI22XLTH U485 ( .A0(n599), .A1(n1745), .B0(n654), .B1(n1747), .Y(n362) );
  OAI22XLTH U486 ( .A0(n599), .A1(n1742), .B0(n653), .B1(n1744), .Y(n363) );
  OAI22XLTH U487 ( .A0(n599), .A1(n1739), .B0(n653), .B1(n1741), .Y(n364) );
  OAI22XLTH U488 ( .A0(n600), .A1(n1736), .B0(n653), .B1(n1738), .Y(n365) );
  OAI22XLTH U489 ( .A0(n600), .A1(n1583), .B0(n653), .B1(n1735), .Y(n366) );
  OAI22XLTH U490 ( .A0(n600), .A1(n1580), .B0(n653), .B1(n1732), .Y(n368) );
  CLKBUFX4TH U491 ( .A(n692), .Y(n691) );
  OAI22XLTH U492 ( .A0(n600), .A1(n1727), .B0(n652), .B1(n1729), .Y(n370) );
  OAI22XLTH U493 ( .A0(n600), .A1(n1724), .B0(n652), .B1(n1726), .Y(n371) );
  CLKBUFX4TH U494 ( .A(n698), .Y(n680) );
  OAI22XLTH U495 ( .A0(n600), .A1(n1721), .B0(n652), .B1(n1723), .Y(n372) );
  OAI22XLTH U496 ( .A0(n600), .A1(n1718), .B0(n651), .B1(n1720), .Y(n373) );
  OAI22XLTH U497 ( .A0(n600), .A1(n1715), .B0(n652), .B1(n1717), .Y(n374) );
  OAI22XLTH U498 ( .A0(n600), .A1(n1712), .B0(n651), .B1(n1714), .Y(n375) );
  OAI22XLTH U499 ( .A0(n600), .A1(n1709), .B0(n651), .B1(n1711), .Y(n376) );
  OAI22XLTH U500 ( .A0(n600), .A1(n1706), .B0(n651), .B1(n1708), .Y(n377) );
  OAI22XLTH U501 ( .A0(n600), .A1(n1703), .B0(n651), .B1(n1705), .Y(n378) );
  OAI22XLTH U502 ( .A0(n601), .A1(n1700), .B0(n650), .B1(n1702), .Y(n379) );
  OAI22XLTH U503 ( .A0(n601), .A1(n2252), .B0(n651), .B1(n1699), .Y(n380) );
  CLKBUFX1TH U504 ( .A(n702), .Y(n701) );
  OAI2B2XLTH U505 ( .A1N(in[2]), .A0(n598), .B0(n2251), .B1(n621), .Y(n381) );
  CLKBUFX4TH U506 ( .A(n699), .Y(n679) );
  OAI2BB2XLTH U507 ( .B0(n598), .B1(n1568), .A0N(n2262), .A1N(n615), .Y(n334)
         );
  OAI2BB1XLTH U508 ( .A0N(N12), .A1N(n654), .B0(n1556), .Y(n486) );
  OAI2BB1XLTH U509 ( .A0N(N11), .A1N(n654), .B0(n1227), .Y(n485) );
  CLKBUFX4TH U510 ( .A(n696), .Y(n685) );
  OAI2BB1XLTH U511 ( .A0N(N13), .A1N(n654), .B0(n1559), .Y(n487) );
  AO22XLTH U512 ( .A0(count2[0]), .A1(n597), .B0(N15), .B1(n1225), .Y(n497) );
  OAI21XLTH U513 ( .A0(n654), .A1(n1562), .B0(n597), .Y(n476) );
  INVXLTH U514 ( .A(out16[0]), .Y(n1294) );
  INVXLTH U515 ( .A(out0[1]), .Y(n1322) );
  INVXLTH U516 ( .A(out45[1]), .Y(n1406) );
  INVXLTH U517 ( .A(out21[1]), .Y(n1384) );
  INVXLTH U518 ( .A(out16[1]), .Y(n1381) );
  INVXLTH U519 ( .A(out45[4]), .Y(n1450) );
  INVXLTH U520 ( .A(out39[4]), .Y(n1444) );
  INVXLTH U521 ( .A(out27[4]), .Y(n1432) );
  INVXLTH U522 ( .A(out16[4]), .Y(n1422) );
  INVXLTH U523 ( .A(out45[2]), .Y(n1366) );
  INVXLTH U524 ( .A(out32[2]), .Y(n1353) );
  INVXLTH U525 ( .A(out46[0]), .Y(n1277) );
  INVXLTH U526 ( .A(out0[0]), .Y(n1278) );
  INVXLTH U527 ( .A(out43[0]), .Y(n1319) );
  INVXLTH U528 ( .A(out42[0]), .Y(n1318) );
  INVXLTH U529 ( .A(out40[0]), .Y(n1316) );
  INVXLTH U530 ( .A(out39[0]), .Y(n1315) );
  INVXLTH U531 ( .A(out38[0]), .Y(n1314) );
  INVXLTH U532 ( .A(out36[0]), .Y(n1312) );
  INVXLTH U533 ( .A(out35[0]), .Y(n1311) );
  INVXLTH U534 ( .A(out33[0]), .Y(n1309) );
  INVXLTH U535 ( .A(out32[0]), .Y(n1308) );
  INVXLTH U536 ( .A(out31[0]), .Y(n1307) );
  INVXLTH U537 ( .A(out30[0]), .Y(n1306) );
  INVXLTH U538 ( .A(out29[0]), .Y(n1305) );
  INVXLTH U539 ( .A(out28[0]), .Y(n1304) );
  INVXLTH U540 ( .A(out27[0]), .Y(n1303) );
  INVXLTH U541 ( .A(out25[0]), .Y(n1301) );
  INVXLTH U542 ( .A(out24[0]), .Y(n1300) );
  INVXLTH U543 ( .A(out22[0]), .Y(n1298) );
  INVXLTH U544 ( .A(out21[0]), .Y(n1297) );
  INVXLTH U545 ( .A(out20[0]), .Y(n1454) );
  INVXLTH U546 ( .A(out19[0]), .Y(n1296) );
  INVXLTH U547 ( .A(out18[0]), .Y(n1295) );
  INVXLTH U548 ( .A(out17[0]), .Y(n1461) );
  INVXLTH U549 ( .A(out15[0]), .Y(n1293) );
  INVXLTH U550 ( .A(out14[0]), .Y(n1292) );
  INVXLTH U551 ( .A(out13[0]), .Y(n1291) );
  INVXLTH U552 ( .A(out12[0]), .Y(n1290) );
  INVXLTH U553 ( .A(out8[0]), .Y(n1286) );
  INVXLTH U554 ( .A(out7[0]), .Y(n1285) );
  INVXLTH U555 ( .A(out6[0]), .Y(n1284) );
  INVXLTH U556 ( .A(out5[0]), .Y(n1283) );
  INVXLTH U557 ( .A(out4[0]), .Y(n1282) );
  INVXLTH U558 ( .A(out1[0]), .Y(n1279) );
  INVXLTH U559 ( .A(out45[0]), .Y(n1276) );
  INVXLTH U560 ( .A(out44[0]), .Y(n1320) );
  INVXLTH U561 ( .A(out3[0]), .Y(n1281) );
  INVXLTH U562 ( .A(out46[1]), .Y(n1407) );
  INVXLTH U563 ( .A(out42[1]), .Y(n1404) );
  INVXLTH U564 ( .A(out39[1]), .Y(n1401) );
  INVXLTH U565 ( .A(out36[1]), .Y(n1399) );
  INVXLTH U566 ( .A(out35[1]), .Y(n1398) );
  INVXLTH U567 ( .A(out33[1]), .Y(n1396) );
  INVXLTH U568 ( .A(out32[1]), .Y(n1395) );
  INVXLTH U569 ( .A(out30[1]), .Y(n1393) );
  INVXLTH U570 ( .A(out29[1]), .Y(n1392) );
  INVXLTH U571 ( .A(out28[1]), .Y(n1391) );
  INVXLTH U572 ( .A(out27[1]), .Y(n1390) );
  INVXLTH U573 ( .A(out24[1]), .Y(n1387) );
  INVXLTH U574 ( .A(out22[1]), .Y(n1385) );
  INVXLTH U575 ( .A(out20[1]), .Y(n1455) );
  INVXLTH U576 ( .A(out19[1]), .Y(n1383) );
  INVXLTH U577 ( .A(out18[1]), .Y(n1382) );
  INVXLTH U578 ( .A(out17[1]), .Y(n1462) );
  INVXLTH U579 ( .A(out15[1]), .Y(n1380) );
  INVXLTH U580 ( .A(out14[1]), .Y(n1379) );
  INVXLTH U581 ( .A(out13[1]), .Y(n1378) );
  INVXLTH U582 ( .A(out12[1]), .Y(n1377) );
  INVXLTH U583 ( .A(out8[1]), .Y(n1374) );
  INVXLTH U584 ( .A(out7[1]), .Y(n1456) );
  INVXLTH U585 ( .A(out4[1]), .Y(n1371) );
  INVXLTH U586 ( .A(out3[1]), .Y(n1370) );
  INVXLTH U587 ( .A(out1[1]), .Y(n1368) );
  INVXLTH U588 ( .A(out36[4]), .Y(n1441) );
  INVXLTH U589 ( .A(out32[4]), .Y(n1437) );
  INVXLTH U590 ( .A(out28[4]), .Y(n1433) );
  INVXLTH U591 ( .A(out20[4]), .Y(n1425) );
  INVXLTH U592 ( .A(out19[4]), .Y(n1424) );
  INVXLTH U593 ( .A(out14[4]), .Y(n1420) );
  INVXLTH U594 ( .A(out13[4]), .Y(n1419) );
  INVXLTH U595 ( .A(out12[4]), .Y(n1418) );
  INVXLTH U596 ( .A(out8[4]), .Y(n1414) );
  INVXLTH U597 ( .A(out4[4]), .Y(n1411) );
  INVXLTH U598 ( .A(out1[4]), .Y(n1408) );
  INVXLTH U599 ( .A(out28[2]), .Y(n1349) );
  INVXLTH U600 ( .A(out14[2]), .Y(n1336) );
  INVXLTH U601 ( .A(out12[2]), .Y(n1334) );
  AOI31XLTH U602 ( .A0(count[5]), .A1(n505), .A2(count[4]), .B0(count[6]), .Y(
        n504) );
  OR4XLTH U603 ( .A(count[3]), .B(count[2]), .C(count[0]), .D(count[1]), .Y(
        n505) );
  OR2XLTH U604 ( .A(count1), .B(n598), .Y(n478) );
  AO22XLTH U605 ( .A0(in[4]), .A1(n617), .B0(n598), .B1(n2263), .Y(n477) );
  AO22XLTH U606 ( .A0(N4), .A1(n619), .B0(n1552), .B1(n599), .Y(n488) );
  AO22XLTH U607 ( .A0(N5), .A1(n617), .B0(count[1]), .B1(n598), .Y(n479) );
  AO22XLTH U608 ( .A0(N6), .A1(n616), .B0(count[2]), .B1(n599), .Y(n480) );
  AO22XLTH U609 ( .A0(N7), .A1(n618), .B0(count[3]), .B1(n598), .Y(n481) );
  AO22XLTH U610 ( .A0(N9), .A1(n616), .B0(count[5]), .B1(n599), .Y(n483) );
  AO22XLTH U611 ( .A0(N8), .A1(n618), .B0(count[4]), .B1(n599), .Y(n482) );
  AO21XLTH U612 ( .A0(N10), .A1(n620), .B0(count[6]), .Y(n484) );
  DLY1X1TH U1133 ( .A(n1507), .Y(n1465) );
  DLY1X1TH U1134 ( .A(n1549), .Y(n1466) );
  DLY1X1TH U1135 ( .A(n1550), .Y(n1467) );
  DLY1X1TH U1136 ( .A(n1520), .Y(n1468) );
  DLY1X1TH U1137 ( .A(n1521), .Y(n1469) );
  DLY1X1TH U1138 ( .A(n1522), .Y(n1470) );
  DLY1X1TH U1139 ( .A(n1523), .Y(n1471) );
  DLY1X1TH U1140 ( .A(n1524), .Y(n1472) );
  DLY1X1TH U1141 ( .A(n1525), .Y(n1473) );
  DLY1X1TH U1142 ( .A(n1526), .Y(n1474) );
  DLY1X1TH U1143 ( .A(n1527), .Y(n1475) );
  DLY1X1TH U1144 ( .A(n1528), .Y(n1476) );
  DLY1X1TH U1145 ( .A(n1529), .Y(n1477) );
  DLY1X1TH U1146 ( .A(n1530), .Y(n1478) );
  DLY1X1TH U1147 ( .A(n1531), .Y(n1479) );
  DLY1X1TH U1148 ( .A(n1532), .Y(n1480) );
  DLY1X1TH U1149 ( .A(n1533), .Y(n1481) );
  DLY1X1TH U1150 ( .A(n1534), .Y(n1482) );
  DLY1X1TH U1151 ( .A(n1535), .Y(n1483) );
  DLY1X1TH U1152 ( .A(n1536), .Y(n1484) );
  DLY1X1TH U1153 ( .A(n1537), .Y(n1485) );
  DLY1X1TH U1154 ( .A(n1538), .Y(n1486) );
  DLY1X1TH U1155 ( .A(n1539), .Y(n1487) );
  DLY1X1TH U1156 ( .A(n1540), .Y(n1488) );
  DLY1X1TH U1157 ( .A(n1541), .Y(n1489) );
  DLY1X1TH U1158 ( .A(n1542), .Y(n1490) );
  DLY1X1TH U1159 ( .A(n1543), .Y(n1491) );
  DLY1X1TH U1160 ( .A(n1544), .Y(n1492) );
  DLY1X1TH U1161 ( .A(n1545), .Y(n1493) );
  DLY1X1TH U1162 ( .A(n1546), .Y(n1494) );
  DLY1X1TH U1163 ( .A(n1547), .Y(n1495) );
  DLY1X1TH U1164 ( .A(n1548), .Y(n1496) );
  DLY1X1TH U1165 ( .A(n1512), .Y(n1497) );
  DLY1X1TH U1166 ( .A(n1513), .Y(n1498) );
  DLY1X1TH U1167 ( .A(n1514), .Y(n1499) );
  DLY1X1TH U1168 ( .A(n1515), .Y(n1500) );
  DLY1X1TH U1169 ( .A(n1516), .Y(n1501) );
  DLY1X1TH U1170 ( .A(n1517), .Y(n1502) );
  DLY1X1TH U1171 ( .A(n1518), .Y(n1503) );
  DLY1X1TH U1172 ( .A(n1519), .Y(n1504) );
  DLY1X1TH U1173 ( .A(n1507), .Y(n1505) );
  DLY1X1TH U1174 ( .A(n1551), .Y(n1506) );
  DLY1X1TH U1175 ( .A(test_se), .Y(n1507) );
  DLY1X1TH U1176 ( .A(n1465), .Y(n1508) );
  DLY1X1TH U1177 ( .A(n1507), .Y(n1509) );
  DLY1X1TH U1178 ( .A(n1507), .Y(n1510) );
  DLY1X1TH U1179 ( .A(n1465), .Y(n1511) );
  DLY1X1TH U1180 ( .A(n1510), .Y(n1512) );
  DLY1X1TH U1181 ( .A(n1497), .Y(n1513) );
  DLY1X1TH U1182 ( .A(n1498), .Y(n1514) );
  DLY1X1TH U1183 ( .A(n1499), .Y(n1515) );
  DLY1X1TH U1184 ( .A(n1500), .Y(n1516) );
  DLY1X1TH U1185 ( .A(n1501), .Y(n1517) );
  DLY1X1TH U1186 ( .A(n1502), .Y(n1518) );
  DLY1X1TH U1187 ( .A(n1503), .Y(n1519) );
  DLY1X1TH U1188 ( .A(n1504), .Y(n1520) );
  DLY1X1TH U1189 ( .A(n1500), .Y(n1521) );
  DLY1X1TH U1190 ( .A(n1469), .Y(n1522) );
  DLY1X1TH U1191 ( .A(n1470), .Y(n1523) );
  DLY1X1TH U1192 ( .A(n1471), .Y(n1524) );
  DLY1X1TH U1193 ( .A(n1472), .Y(n1525) );
  DLY1X1TH U1194 ( .A(n1473), .Y(n1526) );
  DLY1X1TH U1195 ( .A(n1474), .Y(n1527) );
  DLY1X1TH U1196 ( .A(n1475), .Y(n1528) );
  DLY1X1TH U1197 ( .A(n1476), .Y(n1529) );
  DLY1X1TH U1198 ( .A(n1477), .Y(n1530) );
  DLY1X1TH U1199 ( .A(n1478), .Y(n1531) );
  DLY1X1TH U1200 ( .A(n1479), .Y(n1532) );
  DLY1X1TH U1201 ( .A(n1480), .Y(n1533) );
  DLY1X1TH U1202 ( .A(n1481), .Y(n1534) );
  DLY1X1TH U1203 ( .A(n1482), .Y(n1535) );
  DLY1X1TH U1204 ( .A(n1483), .Y(n1536) );
  DLY1X1TH U1205 ( .A(n1484), .Y(n1537) );
  DLY1X1TH U1206 ( .A(n1485), .Y(n1538) );
  DLY1X1TH U1207 ( .A(n1486), .Y(n1539) );
  DLY1X1TH U1208 ( .A(n1487), .Y(n1540) );
  DLY1X1TH U1209 ( .A(n1488), .Y(n1541) );
  DLY1X1TH U1210 ( .A(n1489), .Y(n1542) );
  DLY1X1TH U1211 ( .A(n1490), .Y(n1543) );
  DLY1X1TH U1212 ( .A(n1491), .Y(n1544) );
  DLY1X1TH U1213 ( .A(n1492), .Y(n1545) );
  DLY1X1TH U1214 ( .A(n1493), .Y(n1546) );
  DLY1X1TH U1215 ( .A(n1494), .Y(n1547) );
  DLY1X1TH U1216 ( .A(n1495), .Y(n1548) );
  DLY1X1TH U1217 ( .A(n1473), .Y(n1549) );
  DLY1X1TH U1218 ( .A(n1479), .Y(n1550) );
  DLY1X1TH U1219 ( .A(n1485), .Y(n1551) );
  DLY1X1TH U1220 ( .A(count[0]), .Y(n1552) );
  DLY1X1TH U1221 ( .A(out47[1]), .Y(n1553) );
  INVXLTH U1222 ( .A(n1228), .Y(n1554) );
  INVXLTH U1223 ( .A(n1554), .Y(n1555) );
  INVXLTH U1224 ( .A(n1554), .Y(n1556) );
  INVXLTH U1225 ( .A(n1226), .Y(n1557) );
  INVXLTH U1226 ( .A(n1557), .Y(n1558) );
  INVXLTH U1227 ( .A(n1557), .Y(n1559) );
  INVXLTH U1228 ( .A(n1408), .Y(n1560) );
  INVXLTH U1229 ( .A(n1560), .Y(n1561) );
  INVXLTH U1230 ( .A(n1560), .Y(n1562) );
  INVXLTH U1231 ( .A(n1277), .Y(n1563) );
  INVXLTH U1232 ( .A(n1563), .Y(n1564) );
  INVXLTH U1233 ( .A(n1563), .Y(n1565) );
  INVXLTH U1234 ( .A(n1367), .Y(n1566) );
  INVXLTH U1235 ( .A(n1566), .Y(n1567) );
  INVXLTH U1236 ( .A(n1566), .Y(n1568) );
  INVXLTH U1237 ( .A(n1275), .Y(n1569) );
  INVXLTH U1238 ( .A(n1569), .Y(n1570) );
  INVXLTH U1239 ( .A(n1569), .Y(n1571) );
  INVXLTH U1240 ( .A(n1407), .Y(n1572) );
  INVXLTH U1241 ( .A(n1572), .Y(n1573) );
  INVXLTH U1242 ( .A(n1572), .Y(n1574) );
  INVXLTH U1243 ( .A(n1451), .Y(n1575) );
  INVXLTH U1244 ( .A(n1575), .Y(n1576) );
  INVXLTH U1245 ( .A(n1575), .Y(n1577) );
  INVXLTH U1246 ( .A(n1334), .Y(n1578) );
  INVXLTH U1247 ( .A(n1578), .Y(n1579) );
  INVXLTH U1248 ( .A(n1578), .Y(n1580) );
  INVXLTH U1249 ( .A(n1336), .Y(n1581) );
  INVXLTH U1250 ( .A(n1581), .Y(n1582) );
  INVXLTH U1251 ( .A(n1581), .Y(n1583) );
  INVXLTH U1252 ( .A(n1349), .Y(n1584) );
  INVXLTH U1253 ( .A(n1584), .Y(n1585) );
  INVXLTH U1254 ( .A(n1584), .Y(n1586) );
  INVXLTH U1255 ( .A(n1281), .Y(n1587) );
  INVXLTH U1256 ( .A(n1587), .Y(n1588) );
  INVXLTH U1257 ( .A(n1587), .Y(n1589) );
  INVXLTH U1258 ( .A(n1320), .Y(n1590) );
  INVXLTH U1259 ( .A(n1590), .Y(n1591) );
  INVXLTH U1260 ( .A(n1590), .Y(n1592) );
  INVXLTH U1261 ( .A(n1276), .Y(n1593) );
  INVXLTH U1262 ( .A(n1593), .Y(n1594) );
  INVXLTH U1263 ( .A(n1593), .Y(n1595) );
  INVXLTH U1264 ( .A(n1279), .Y(n1596) );
  INVXLTH U1265 ( .A(n1596), .Y(n1597) );
  INVXLTH U1266 ( .A(n1596), .Y(n1598) );
  INVXLTH U1267 ( .A(n1282), .Y(n1599) );
  INVXLTH U1268 ( .A(n1599), .Y(n1600) );
  INVXLTH U1269 ( .A(n1599), .Y(n1601) );
  INVXLTH U1270 ( .A(n1283), .Y(n1602) );
  INVXLTH U1271 ( .A(n1602), .Y(n1603) );
  INVXLTH U1272 ( .A(n1602), .Y(n1604) );
  INVXLTH U1273 ( .A(n1284), .Y(n1605) );
  INVXLTH U1274 ( .A(n1605), .Y(n1606) );
  INVXLTH U1275 ( .A(n1605), .Y(n1607) );
  INVXLTH U1276 ( .A(n1285), .Y(n1608) );
  INVXLTH U1277 ( .A(n1608), .Y(n1609) );
  INVXLTH U1278 ( .A(n1608), .Y(n1610) );
  INVXLTH U1279 ( .A(n1286), .Y(n1611) );
  INVXLTH U1280 ( .A(n1611), .Y(n1612) );
  INVXLTH U1281 ( .A(n1611), .Y(n1613) );
  INVXLTH U1282 ( .A(n1290), .Y(n1614) );
  INVXLTH U1283 ( .A(n1614), .Y(n1615) );
  INVXLTH U1284 ( .A(n1614), .Y(n1616) );
  INVXLTH U1285 ( .A(n1291), .Y(n1617) );
  INVXLTH U1286 ( .A(n1617), .Y(n1618) );
  INVXLTH U1287 ( .A(n1617), .Y(n1619) );
  INVXLTH U1288 ( .A(n1292), .Y(n1620) );
  INVXLTH U1289 ( .A(n1620), .Y(n1621) );
  INVXLTH U1290 ( .A(n1620), .Y(n1622) );
  INVXLTH U1291 ( .A(n1293), .Y(n1623) );
  INVXLTH U1292 ( .A(n1623), .Y(n1624) );
  INVXLTH U1293 ( .A(n1623), .Y(n1625) );
  INVXLTH U1294 ( .A(n1461), .Y(n1626) );
  INVXLTH U1295 ( .A(n1626), .Y(n1627) );
  INVXLTH U1296 ( .A(n1626), .Y(n1628) );
  INVXLTH U1297 ( .A(n1295), .Y(n1629) );
  INVXLTH U1298 ( .A(n1629), .Y(n1630) );
  INVXLTH U1299 ( .A(n1629), .Y(n1631) );
  INVXLTH U1300 ( .A(n1296), .Y(n1632) );
  INVXLTH U1301 ( .A(n1632), .Y(n1633) );
  INVXLTH U1302 ( .A(n1632), .Y(n1634) );
  INVXLTH U1303 ( .A(n1454), .Y(n1635) );
  INVXLTH U1304 ( .A(n1635), .Y(n1636) );
  INVXLTH U1305 ( .A(n1635), .Y(n1637) );
  INVXLTH U1306 ( .A(n1297), .Y(n1638) );
  INVXLTH U1307 ( .A(n1638), .Y(n1639) );
  INVXLTH U1308 ( .A(n1638), .Y(n1640) );
  INVXLTH U1309 ( .A(n1298), .Y(n1641) );
  INVXLTH U1310 ( .A(n1641), .Y(n1642) );
  INVXLTH U1311 ( .A(n1641), .Y(n1643) );
  INVXLTH U1312 ( .A(n1300), .Y(n1644) );
  INVXLTH U1313 ( .A(n1644), .Y(n1645) );
  INVXLTH U1314 ( .A(n1644), .Y(n1646) );
  INVXLTH U1315 ( .A(n1301), .Y(n1647) );
  INVXLTH U1316 ( .A(n1647), .Y(n1648) );
  INVXLTH U1317 ( .A(n1647), .Y(n1649) );
  INVXLTH U1318 ( .A(n1303), .Y(n1650) );
  INVXLTH U1319 ( .A(n1650), .Y(n1651) );
  INVXLTH U1320 ( .A(n1650), .Y(n1652) );
  INVXLTH U1321 ( .A(n1304), .Y(n1653) );
  INVXLTH U1322 ( .A(n1653), .Y(n1654) );
  INVXLTH U1323 ( .A(n1653), .Y(n1655) );
  INVXLTH U1324 ( .A(n1305), .Y(n1656) );
  INVXLTH U1325 ( .A(n1656), .Y(n1657) );
  INVXLTH U1326 ( .A(n1656), .Y(n1658) );
  INVXLTH U1327 ( .A(n1306), .Y(n1659) );
  INVXLTH U1328 ( .A(n1659), .Y(n1660) );
  INVXLTH U1329 ( .A(n1659), .Y(n1661) );
  INVXLTH U1330 ( .A(n1307), .Y(n1662) );
  INVXLTH U1331 ( .A(n1662), .Y(n1663) );
  INVXLTH U1332 ( .A(n1662), .Y(n1664) );
  INVXLTH U1333 ( .A(n1308), .Y(n1665) );
  INVXLTH U1334 ( .A(n1665), .Y(n1666) );
  INVXLTH U1335 ( .A(n1665), .Y(n1667) );
  INVXLTH U1336 ( .A(n1309), .Y(n1668) );
  INVXLTH U1337 ( .A(n1668), .Y(n1669) );
  INVXLTH U1338 ( .A(n1668), .Y(n1670) );
  INVXLTH U1339 ( .A(n1311), .Y(n1671) );
  INVXLTH U1340 ( .A(n1671), .Y(n1672) );
  INVXLTH U1341 ( .A(n1671), .Y(n1673) );
  INVXLTH U1342 ( .A(n1312), .Y(n1674) );
  INVXLTH U1343 ( .A(n1674), .Y(n1675) );
  INVXLTH U1344 ( .A(n1674), .Y(n1676) );
  INVXLTH U1345 ( .A(n1314), .Y(n1677) );
  INVXLTH U1346 ( .A(n1677), .Y(n1678) );
  INVXLTH U1347 ( .A(n1677), .Y(n1679) );
  INVXLTH U1348 ( .A(n1315), .Y(n1680) );
  INVXLTH U1349 ( .A(n1680), .Y(n1681) );
  INVXLTH U1350 ( .A(n1680), .Y(n1682) );
  INVXLTH U1351 ( .A(n1316), .Y(n1683) );
  INVXLTH U1352 ( .A(n1683), .Y(n1684) );
  INVXLTH U1353 ( .A(n1683), .Y(n1685) );
  INVXLTH U1354 ( .A(n1319), .Y(n1686) );
  INVXLTH U1355 ( .A(n1686), .Y(n1687) );
  INVXLTH U1356 ( .A(n1686), .Y(n1688) );
  INVXLTH U1357 ( .A(n1353), .Y(n1689) );
  INVXLTH U1358 ( .A(n1689), .Y(n1690) );
  INVXLTH U1359 ( .A(n1689), .Y(n1691) );
  INVXLTH U1360 ( .A(n1366), .Y(n1692) );
  INVXLTH U1361 ( .A(n1692), .Y(n1693) );
  INVXLTH U1362 ( .A(n1692), .Y(n1694) );
  INVXLTH U1363 ( .A(n1294), .Y(n1695) );
  INVXLTH U1364 ( .A(n1695), .Y(n1696) );
  INVXLTH U1365 ( .A(n1695), .Y(n1697) );
  INVXLTH U1366 ( .A(n1323), .Y(n1698) );
  INVXLTH U1367 ( .A(n1698), .Y(n1699) );
  INVXLTH U1368 ( .A(n1698), .Y(n1700) );
  INVXLTH U1369 ( .A(n1324), .Y(n1701) );
  INVXLTH U1370 ( .A(n1701), .Y(n1702) );
  INVXLTH U1371 ( .A(n1701), .Y(n1703) );
  INVXLTH U1372 ( .A(n1325), .Y(n1704) );
  INVXLTH U1373 ( .A(n1704), .Y(n1705) );
  INVXLTH U1374 ( .A(n1704), .Y(n1706) );
  INVXLTH U1375 ( .A(n1326), .Y(n1707) );
  INVXLTH U1376 ( .A(n1707), .Y(n1708) );
  INVXLTH U1377 ( .A(n1707), .Y(n1709) );
  INVXLTH U1378 ( .A(n1327), .Y(n1710) );
  INVXLTH U1379 ( .A(n1710), .Y(n1711) );
  INVXLTH U1380 ( .A(n1710), .Y(n1712) );
  INVXLTH U1381 ( .A(n1328), .Y(n1713) );
  INVXLTH U1382 ( .A(n1713), .Y(n1714) );
  INVXLTH U1383 ( .A(n1713), .Y(n1715) );
  INVXLTH U1384 ( .A(n1329), .Y(n1716) );
  INVXLTH U1385 ( .A(n1716), .Y(n1717) );
  INVXLTH U1386 ( .A(n1716), .Y(n1718) );
  INVXLTH U1387 ( .A(n1330), .Y(n1719) );
  INVXLTH U1388 ( .A(n1719), .Y(n1720) );
  INVXLTH U1389 ( .A(n1719), .Y(n1721) );
  INVXLTH U1390 ( .A(n1331), .Y(n1722) );
  INVXLTH U1391 ( .A(n1722), .Y(n1723) );
  INVXLTH U1392 ( .A(n1722), .Y(n1724) );
  INVXLTH U1393 ( .A(n1332), .Y(n1725) );
  INVXLTH U1394 ( .A(n1725), .Y(n1726) );
  INVXLTH U1395 ( .A(n1725), .Y(n1727) );
  INVXLTH U1396 ( .A(n1333), .Y(n1728) );
  INVXLTH U1397 ( .A(n1728), .Y(n1729) );
  INVXLTH U1398 ( .A(n1728), .Y(n1730) );
  INVXLTH U1399 ( .A(n1335), .Y(n1731) );
  INVXLTH U1400 ( .A(n1731), .Y(n1732) );
  INVXLTH U1401 ( .A(n1731), .Y(n1733) );
  INVXLTH U1402 ( .A(n1337), .Y(n1734) );
  INVXLTH U1403 ( .A(n1734), .Y(n1735) );
  INVXLTH U1404 ( .A(n1734), .Y(n1736) );
  INVXLTH U1405 ( .A(n1338), .Y(n1737) );
  INVXLTH U1406 ( .A(n1737), .Y(n1738) );
  INVXLTH U1407 ( .A(n1737), .Y(n1739) );
  INVXLTH U1408 ( .A(n1339), .Y(n1740) );
  INVXLTH U1409 ( .A(n1740), .Y(n1741) );
  INVXLTH U1410 ( .A(n1740), .Y(n1742) );
  INVXLTH U1411 ( .A(n1340), .Y(n1743) );
  INVXLTH U1412 ( .A(n1743), .Y(n1744) );
  INVXLTH U1413 ( .A(n1743), .Y(n1745) );
  INVXLTH U1414 ( .A(n1341), .Y(n1746) );
  INVXLTH U1415 ( .A(n1746), .Y(n1747) );
  INVXLTH U1416 ( .A(n1746), .Y(n1748) );
  INVXLTH U1417 ( .A(n1342), .Y(n1749) );
  INVXLTH U1418 ( .A(n1749), .Y(n1750) );
  INVXLTH U1419 ( .A(n1749), .Y(n1751) );
  INVXLTH U1420 ( .A(n1343), .Y(n1752) );
  INVXLTH U1421 ( .A(n1752), .Y(n1753) );
  INVXLTH U1422 ( .A(n1752), .Y(n1754) );
  INVXLTH U1423 ( .A(n1344), .Y(n1755) );
  INVXLTH U1424 ( .A(n1755), .Y(n1756) );
  INVXLTH U1425 ( .A(n1755), .Y(n1757) );
  INVXLTH U1426 ( .A(n1345), .Y(n1758) );
  INVXLTH U1427 ( .A(n1758), .Y(n1759) );
  INVXLTH U1428 ( .A(n1758), .Y(n1760) );
  INVXLTH U1429 ( .A(n1346), .Y(n1761) );
  INVXLTH U1430 ( .A(n1761), .Y(n1762) );
  INVXLTH U1431 ( .A(n1761), .Y(n1763) );
  INVXLTH U1432 ( .A(n1347), .Y(n1764) );
  INVXLTH U1433 ( .A(n1764), .Y(n1765) );
  INVXLTH U1434 ( .A(n1764), .Y(n1766) );
  INVXLTH U1435 ( .A(n1460), .Y(n1767) );
  INVXLTH U1436 ( .A(n1767), .Y(n1768) );
  INVXLTH U1437 ( .A(n1767), .Y(n1769) );
  INVXLTH U1438 ( .A(n1348), .Y(n1770) );
  INVXLTH U1439 ( .A(n1770), .Y(n1771) );
  INVXLTH U1440 ( .A(n1770), .Y(n1772) );
  INVXLTH U1441 ( .A(n1350), .Y(n1773) );
  INVXLTH U1442 ( .A(n1773), .Y(n1774) );
  INVXLTH U1443 ( .A(n1773), .Y(n1775) );
  INVXLTH U1444 ( .A(n1351), .Y(n1776) );
  INVXLTH U1445 ( .A(n1776), .Y(n1777) );
  INVXLTH U1446 ( .A(n1776), .Y(n1778) );
  INVXLTH U1447 ( .A(n1352), .Y(n1779) );
  INVXLTH U1448 ( .A(n1779), .Y(n1780) );
  INVXLTH U1449 ( .A(n1779), .Y(n1781) );
  INVXLTH U1450 ( .A(n1354), .Y(n1782) );
  INVXLTH U1451 ( .A(n1782), .Y(n1783) );
  INVXLTH U1452 ( .A(n1782), .Y(n1784) );
  INVXLTH U1453 ( .A(n1355), .Y(n1785) );
  INVXLTH U1454 ( .A(n1785), .Y(n1786) );
  INVXLTH U1455 ( .A(n1785), .Y(n1787) );
  INVXLTH U1456 ( .A(n1356), .Y(n1788) );
  INVXLTH U1457 ( .A(n1788), .Y(n1789) );
  INVXLTH U1458 ( .A(n1788), .Y(n1790) );
  INVXLTH U1459 ( .A(n1357), .Y(n1791) );
  INVXLTH U1460 ( .A(n1791), .Y(n1792) );
  INVXLTH U1461 ( .A(n1791), .Y(n1793) );
  INVXLTH U1462 ( .A(n1358), .Y(n1794) );
  INVXLTH U1463 ( .A(n1794), .Y(n1795) );
  INVXLTH U1464 ( .A(n1794), .Y(n1796) );
  INVXLTH U1465 ( .A(n1359), .Y(n1797) );
  INVXLTH U1466 ( .A(n1797), .Y(n1798) );
  INVXLTH U1467 ( .A(n1797), .Y(n1799) );
  INVXLTH U1468 ( .A(n1360), .Y(n1800) );
  INVXLTH U1469 ( .A(n1800), .Y(n1801) );
  INVXLTH U1470 ( .A(n1800), .Y(n1802) );
  INVXLTH U1471 ( .A(n1361), .Y(n1803) );
  INVXLTH U1472 ( .A(n1803), .Y(n1804) );
  INVXLTH U1473 ( .A(n1803), .Y(n1805) );
  INVXLTH U1474 ( .A(n1362), .Y(n1806) );
  INVXLTH U1475 ( .A(n1806), .Y(n1807) );
  INVXLTH U1476 ( .A(n1806), .Y(n1808) );
  INVXLTH U1477 ( .A(n1363), .Y(n1809) );
  INVXLTH U1478 ( .A(n1809), .Y(n1810) );
  INVXLTH U1479 ( .A(n1809), .Y(n1811) );
  INVXLTH U1480 ( .A(n1364), .Y(n1812) );
  INVXLTH U1481 ( .A(n1812), .Y(n1813) );
  INVXLTH U1482 ( .A(n1812), .Y(n1814) );
  INVXLTH U1483 ( .A(n1365), .Y(n1815) );
  INVXLTH U1484 ( .A(n1815), .Y(n1816) );
  INVXLTH U1485 ( .A(n1815), .Y(n1817) );
  INVXLTH U1486 ( .A(n1302), .Y(n1818) );
  INVXLTH U1487 ( .A(n1818), .Y(n1819) );
  INVXLTH U1488 ( .A(n1818), .Y(n1820) );
  INVXLTH U1489 ( .A(n1280), .Y(n1821) );
  INVXLTH U1490 ( .A(n1821), .Y(n1822) );
  INVXLTH U1491 ( .A(n1821), .Y(n1823) );
  INVXLTH U1492 ( .A(n1313), .Y(n1824) );
  INVXLTH U1493 ( .A(n1824), .Y(n1825) );
  INVXLTH U1494 ( .A(n1824), .Y(n1826) );
  INVXLTH U1495 ( .A(n1317), .Y(n1827) );
  INVXLTH U1496 ( .A(n1827), .Y(n1828) );
  INVXLTH U1497 ( .A(n1827), .Y(n1829) );
  INVXLTH U1498 ( .A(n1299), .Y(n1830) );
  INVXLTH U1499 ( .A(n1830), .Y(n1831) );
  INVXLTH U1500 ( .A(n1830), .Y(n1832) );
  INVXLTH U1501 ( .A(n1310), .Y(n1833) );
  INVXLTH U1502 ( .A(n1833), .Y(n1834) );
  INVXLTH U1503 ( .A(n1833), .Y(n1835) );
  INVXLTH U1504 ( .A(n1289), .Y(n1836) );
  INVXLTH U1505 ( .A(n1836), .Y(n1837) );
  INVXLTH U1506 ( .A(n1836), .Y(n1838) );
  INVXLTH U1507 ( .A(n1242), .Y(n1839) );
  INVXLTH U1508 ( .A(n1839), .Y(n1840) );
  INVXLTH U1509 ( .A(n1839), .Y(n1841) );
  INVXLTH U1510 ( .A(n1243), .Y(n1842) );
  INVXLTH U1511 ( .A(n1842), .Y(n1843) );
  INVXLTH U1512 ( .A(n1842), .Y(n1844) );
  INVXLTH U1513 ( .A(n1232), .Y(n1845) );
  INVXLTH U1514 ( .A(n1845), .Y(n1846) );
  INVXLTH U1515 ( .A(n1845), .Y(n1847) );
  INVXLTH U1516 ( .A(n1233), .Y(n1848) );
  INVXLTH U1517 ( .A(n1848), .Y(n1849) );
  INVXLTH U1518 ( .A(n1848), .Y(n1850) );
  INVXLTH U1519 ( .A(n1247), .Y(n1851) );
  INVXLTH U1520 ( .A(n1851), .Y(n1852) );
  INVXLTH U1521 ( .A(n1851), .Y(n1853) );
  INVXLTH U1522 ( .A(n1248), .Y(n1854) );
  INVXLTH U1523 ( .A(n1854), .Y(n1855) );
  INVXLTH U1524 ( .A(n1854), .Y(n1856) );
  INVXLTH U1525 ( .A(n1249), .Y(n1857) );
  INVXLTH U1526 ( .A(n1857), .Y(n1858) );
  INVXLTH U1527 ( .A(n1857), .Y(n1859) );
  INVXLTH U1528 ( .A(n1256), .Y(n1860) );
  INVXLTH U1529 ( .A(n1860), .Y(n1861) );
  INVXLTH U1530 ( .A(n1860), .Y(n1862) );
  INVXLTH U1531 ( .A(n1257), .Y(n1863) );
  INVXLTH U1532 ( .A(n1863), .Y(n1864) );
  INVXLTH U1533 ( .A(n1863), .Y(n1865) );
  INVXLTH U1534 ( .A(n1265), .Y(n1866) );
  INVXLTH U1535 ( .A(n1866), .Y(n1867) );
  INVXLTH U1536 ( .A(n1866), .Y(n1868) );
  INVXLTH U1537 ( .A(n1264), .Y(n1869) );
  INVXLTH U1538 ( .A(n1869), .Y(n1870) );
  INVXLTH U1539 ( .A(n1869), .Y(n1871) );
  INVXLTH U1540 ( .A(n1231), .Y(n1872) );
  INVXLTH U1541 ( .A(n1872), .Y(n1873) );
  INVXLTH U1542 ( .A(n1872), .Y(n1874) );
  INVXLTH U1543 ( .A(n1234), .Y(n1875) );
  INVXLTH U1544 ( .A(n1875), .Y(n1876) );
  INVXLTH U1545 ( .A(n1875), .Y(n1877) );
  INVXLTH U1546 ( .A(n1235), .Y(n1878) );
  INVXLTH U1547 ( .A(n1878), .Y(n1879) );
  INVXLTH U1548 ( .A(n1878), .Y(n1880) );
  INVXLTH U1549 ( .A(n1244), .Y(n1881) );
  INVXLTH U1550 ( .A(n1881), .Y(n1882) );
  INVXLTH U1551 ( .A(n1881), .Y(n1883) );
  INVXLTH U1552 ( .A(n1246), .Y(n1884) );
  INVXLTH U1553 ( .A(n1884), .Y(n1885) );
  INVXLTH U1554 ( .A(n1884), .Y(n1886) );
  INVXLTH U1555 ( .A(n1250), .Y(n1887) );
  INVXLTH U1556 ( .A(n1887), .Y(n1888) );
  INVXLTH U1557 ( .A(n1887), .Y(n1889) );
  INVXLTH U1558 ( .A(n1251), .Y(n1890) );
  INVXLTH U1559 ( .A(n1890), .Y(n1891) );
  INVXLTH U1560 ( .A(n1890), .Y(n1892) );
  INVXLTH U1561 ( .A(n1253), .Y(n1893) );
  INVXLTH U1562 ( .A(n1893), .Y(n1894) );
  INVXLTH U1563 ( .A(n1893), .Y(n1895) );
  INVXLTH U1564 ( .A(n1252), .Y(n1896) );
  INVXLTH U1565 ( .A(n1896), .Y(n1897) );
  INVXLTH U1566 ( .A(n1896), .Y(n1898) );
  INVXLTH U1567 ( .A(n1254), .Y(n1899) );
  INVXLTH U1568 ( .A(n1899), .Y(n1900) );
  INVXLTH U1569 ( .A(n1899), .Y(n1901) );
  INVXLTH U1570 ( .A(n1255), .Y(n1902) );
  INVXLTH U1571 ( .A(n1902), .Y(n1903) );
  INVXLTH U1572 ( .A(n1902), .Y(n1904) );
  INVXLTH U1573 ( .A(n1259), .Y(n1905) );
  INVXLTH U1574 ( .A(n1905), .Y(n1906) );
  INVXLTH U1575 ( .A(n1905), .Y(n1907) );
  INVXLTH U1576 ( .A(n1258), .Y(n1908) );
  INVXLTH U1577 ( .A(n1908), .Y(n1909) );
  INVXLTH U1578 ( .A(n1908), .Y(n1910) );
  INVXLTH U1579 ( .A(n1260), .Y(n1911) );
  INVXLTH U1580 ( .A(n1911), .Y(n1912) );
  INVXLTH U1581 ( .A(n1911), .Y(n1913) );
  INVXLTH U1582 ( .A(n1263), .Y(n1914) );
  INVXLTH U1583 ( .A(n1914), .Y(n1915) );
  INVXLTH U1584 ( .A(n1914), .Y(n1916) );
  INVXLTH U1585 ( .A(n1266), .Y(n1917) );
  INVXLTH U1586 ( .A(n1917), .Y(n1918) );
  INVXLTH U1587 ( .A(n1917), .Y(n1919) );
  INVXLTH U1588 ( .A(n1267), .Y(n1920) );
  INVXLTH U1589 ( .A(n1920), .Y(n1921) );
  INVXLTH U1590 ( .A(n1920), .Y(n1922) );
  INVXLTH U1591 ( .A(n1268), .Y(n1923) );
  INVXLTH U1592 ( .A(n1923), .Y(n1924) );
  INVXLTH U1593 ( .A(n1923), .Y(n1925) );
  INVXLTH U1594 ( .A(n1269), .Y(n1926) );
  INVXLTH U1595 ( .A(n1926), .Y(n1927) );
  INVXLTH U1596 ( .A(n1926), .Y(n1928) );
  INVXLTH U1597 ( .A(n1270), .Y(n1929) );
  INVXLTH U1598 ( .A(n1929), .Y(n1930) );
  INVXLTH U1599 ( .A(n1929), .Y(n1931) );
  INVXLTH U1600 ( .A(n1271), .Y(n1932) );
  INVXLTH U1601 ( .A(n1932), .Y(n1933) );
  INVXLTH U1602 ( .A(n1932), .Y(n1934) );
  INVXLTH U1603 ( .A(n1272), .Y(n1935) );
  INVXLTH U1604 ( .A(n1935), .Y(n1936) );
  INVXLTH U1605 ( .A(n1935), .Y(n1937) );
  INVXLTH U1606 ( .A(n1273), .Y(n1938) );
  INVXLTH U1607 ( .A(n1938), .Y(n1939) );
  INVXLTH U1608 ( .A(n1938), .Y(n1940) );
  INVXLTH U1609 ( .A(n1274), .Y(n1941) );
  INVXLTH U1610 ( .A(n1941), .Y(n1942) );
  INVXLTH U1611 ( .A(n1941), .Y(n1943) );
  INVXLTH U1612 ( .A(n1230), .Y(n1944) );
  INVXLTH U1613 ( .A(n1944), .Y(n1945) );
  INVXLTH U1614 ( .A(n1944), .Y(n1946) );
  INVXLTH U1615 ( .A(n1237), .Y(n1947) );
  INVXLTH U1616 ( .A(n1947), .Y(n1948) );
  INVXLTH U1617 ( .A(n1947), .Y(n1949) );
  INVXLTH U1618 ( .A(n1238), .Y(n1950) );
  INVXLTH U1619 ( .A(n1950), .Y(n1951) );
  INVXLTH U1620 ( .A(n1950), .Y(n1952) );
  INVXLTH U1621 ( .A(n1239), .Y(n1953) );
  INVXLTH U1622 ( .A(n1953), .Y(n1954) );
  INVXLTH U1623 ( .A(n1953), .Y(n1955) );
  INVXLTH U1624 ( .A(n1240), .Y(n1956) );
  INVXLTH U1625 ( .A(n1956), .Y(n1957) );
  INVXLTH U1626 ( .A(n1956), .Y(n1958) );
  INVXLTH U1627 ( .A(n1245), .Y(n1959) );
  INVXLTH U1628 ( .A(n1959), .Y(n1960) );
  INVXLTH U1629 ( .A(n1959), .Y(n1961) );
  INVXLTH U1630 ( .A(n1261), .Y(n1962) );
  INVXLTH U1631 ( .A(n1962), .Y(n1963) );
  INVXLTH U1632 ( .A(n1962), .Y(n1964) );
  INVXLTH U1633 ( .A(n1262), .Y(n1965) );
  INVXLTH U1634 ( .A(n1965), .Y(n1966) );
  INVXLTH U1635 ( .A(n1965), .Y(n1967) );
  INVXLTH U1636 ( .A(n1241), .Y(n1968) );
  INVXLTH U1637 ( .A(n1968), .Y(n1969) );
  INVXLTH U1638 ( .A(n1968), .Y(n1970) );
  INVXLTH U1639 ( .A(n1287), .Y(n1971) );
  INVXLTH U1640 ( .A(n1971), .Y(n1972) );
  INVXLTH U1641 ( .A(n1971), .Y(n1973) );
  INVXLTH U1642 ( .A(n1288), .Y(n1974) );
  INVXLTH U1643 ( .A(n1974), .Y(n1975) );
  INVXLTH U1644 ( .A(n1974), .Y(n1976) );
  INVXLTH U1645 ( .A(n1458), .Y(n1977) );
  INVXLTH U1646 ( .A(n1977), .Y(n1978) );
  INVXLTH U1647 ( .A(n1977), .Y(n1979) );
  INVXLTH U1648 ( .A(n1411), .Y(n1980) );
  INVXLTH U1649 ( .A(n1980), .Y(n1981) );
  INVXLTH U1650 ( .A(n1980), .Y(n1982) );
  INVXLTH U1651 ( .A(n1414), .Y(n1983) );
  INVXLTH U1652 ( .A(n1983), .Y(n1984) );
  INVXLTH U1653 ( .A(n1983), .Y(n1985) );
  INVXLTH U1654 ( .A(n1418), .Y(n1986) );
  INVXLTH U1655 ( .A(n1986), .Y(n1987) );
  INVXLTH U1656 ( .A(n1986), .Y(n1988) );
  INVXLTH U1657 ( .A(n1419), .Y(n1989) );
  INVXLTH U1658 ( .A(n1989), .Y(n1990) );
  INVXLTH U1659 ( .A(n1989), .Y(n1991) );
  INVXLTH U1660 ( .A(n1420), .Y(n1992) );
  INVXLTH U1661 ( .A(n1992), .Y(n1993) );
  INVXLTH U1662 ( .A(n1992), .Y(n1994) );
  INVXLTH U1663 ( .A(n1424), .Y(n1995) );
  INVXLTH U1664 ( .A(n1995), .Y(n1996) );
  INVXLTH U1665 ( .A(n1995), .Y(n1997) );
  INVXLTH U1666 ( .A(n1425), .Y(n1998) );
  INVXLTH U1667 ( .A(n1998), .Y(n1999) );
  INVXLTH U1668 ( .A(n1998), .Y(n2000) );
  INVXLTH U1669 ( .A(n1433), .Y(n2001) );
  INVXLTH U1670 ( .A(n2001), .Y(n2002) );
  INVXLTH U1671 ( .A(n2001), .Y(n2003) );
  INVXLTH U1672 ( .A(n1437), .Y(n2004) );
  INVXLTH U1673 ( .A(n2004), .Y(n2005) );
  INVXLTH U1674 ( .A(n2004), .Y(n2006) );
  INVXLTH U1675 ( .A(n1441), .Y(n2007) );
  INVXLTH U1676 ( .A(n2007), .Y(n2008) );
  INVXLTH U1677 ( .A(n2007), .Y(n2009) );
  INVXLTH U1678 ( .A(n1368), .Y(n2010) );
  INVXLTH U1679 ( .A(n2010), .Y(n2011) );
  INVXLTH U1680 ( .A(n2010), .Y(n2012) );
  INVXLTH U1681 ( .A(n1370), .Y(n2013) );
  INVXLTH U1682 ( .A(n2013), .Y(n2014) );
  INVXLTH U1683 ( .A(n2013), .Y(n2015) );
  INVXLTH U1684 ( .A(n1371), .Y(n2016) );
  INVXLTH U1685 ( .A(n2016), .Y(n2017) );
  INVXLTH U1686 ( .A(n2016), .Y(n2018) );
  INVXLTH U1687 ( .A(n1456), .Y(n2019) );
  INVXLTH U1688 ( .A(n2019), .Y(n2020) );
  INVXLTH U1689 ( .A(n2019), .Y(n2021) );
  INVXLTH U1690 ( .A(n1374), .Y(n2022) );
  INVXLTH U1691 ( .A(n2022), .Y(n2023) );
  INVXLTH U1692 ( .A(n2022), .Y(n2024) );
  INVXLTH U1693 ( .A(n1377), .Y(n2025) );
  INVXLTH U1694 ( .A(n2025), .Y(n2026) );
  INVXLTH U1695 ( .A(n2025), .Y(n2027) );
  INVXLTH U1696 ( .A(n1378), .Y(n2028) );
  INVXLTH U1697 ( .A(n2028), .Y(n2029) );
  INVXLTH U1698 ( .A(n2028), .Y(n2030) );
  INVXLTH U1699 ( .A(n1379), .Y(n2031) );
  INVXLTH U1700 ( .A(n2031), .Y(n2032) );
  INVXLTH U1701 ( .A(n2031), .Y(n2033) );
  INVXLTH U1702 ( .A(n1380), .Y(n2034) );
  INVXLTH U1703 ( .A(n2034), .Y(n2035) );
  INVXLTH U1704 ( .A(n2034), .Y(n2036) );
  INVXLTH U1705 ( .A(n1462), .Y(n2037) );
  INVXLTH U1706 ( .A(n2037), .Y(n2038) );
  INVXLTH U1707 ( .A(n2037), .Y(n2039) );
  INVXLTH U1708 ( .A(n1382), .Y(n2040) );
  INVXLTH U1709 ( .A(n2040), .Y(n2041) );
  INVXLTH U1710 ( .A(n2040), .Y(n2042) );
  INVXLTH U1711 ( .A(n1383), .Y(n2043) );
  INVXLTH U1712 ( .A(n2043), .Y(n2044) );
  INVXLTH U1713 ( .A(n2043), .Y(n2045) );
  INVXLTH U1714 ( .A(n1455), .Y(n2046) );
  INVXLTH U1715 ( .A(n2046), .Y(n2047) );
  INVXLTH U1716 ( .A(n2046), .Y(n2048) );
  INVXLTH U1717 ( .A(n1385), .Y(n2049) );
  INVXLTH U1718 ( .A(n2049), .Y(n2050) );
  INVXLTH U1719 ( .A(n2049), .Y(n2051) );
  INVXLTH U1720 ( .A(n1387), .Y(n2052) );
  INVXLTH U1721 ( .A(n2052), .Y(n2053) );
  INVXLTH U1722 ( .A(n2052), .Y(n2054) );
  INVXLTH U1723 ( .A(n1390), .Y(n2055) );
  INVXLTH U1724 ( .A(n2055), .Y(n2056) );
  INVXLTH U1725 ( .A(n2055), .Y(n2057) );
  INVXLTH U1726 ( .A(n1391), .Y(n2058) );
  INVXLTH U1727 ( .A(n2058), .Y(n2059) );
  INVXLTH U1728 ( .A(n2058), .Y(n2060) );
  INVXLTH U1729 ( .A(n1392), .Y(n2061) );
  INVXLTH U1730 ( .A(n2061), .Y(n2062) );
  INVXLTH U1731 ( .A(n2061), .Y(n2063) );
  INVXLTH U1732 ( .A(n1393), .Y(n2064) );
  INVXLTH U1733 ( .A(n2064), .Y(n2065) );
  INVXLTH U1734 ( .A(n2064), .Y(n2066) );
  INVXLTH U1735 ( .A(n1395), .Y(n2067) );
  INVXLTH U1736 ( .A(n2067), .Y(n2068) );
  INVXLTH U1737 ( .A(n2067), .Y(n2069) );
  INVXLTH U1738 ( .A(n1396), .Y(n2070) );
  INVXLTH U1739 ( .A(n2070), .Y(n2071) );
  INVXLTH U1740 ( .A(n2070), .Y(n2072) );
  INVXLTH U1741 ( .A(n1398), .Y(n2073) );
  INVXLTH U1742 ( .A(n2073), .Y(n2074) );
  INVXLTH U1743 ( .A(n2073), .Y(n2075) );
  INVXLTH U1744 ( .A(n1399), .Y(n2076) );
  INVXLTH U1745 ( .A(n2076), .Y(n2077) );
  INVXLTH U1746 ( .A(n2076), .Y(n2078) );
  INVXLTH U1747 ( .A(n1401), .Y(n2079) );
  INVXLTH U1748 ( .A(n2079), .Y(n2080) );
  INVXLTH U1749 ( .A(n2079), .Y(n2081) );
  INVXLTH U1750 ( .A(n1404), .Y(n2082) );
  INVXLTH U1751 ( .A(n2082), .Y(n2083) );
  INVXLTH U1752 ( .A(n2082), .Y(n2084) );
  INVXLTH U1753 ( .A(n1318), .Y(n2085) );
  INVXLTH U1754 ( .A(n2085), .Y(n2086) );
  INVXLTH U1755 ( .A(n2085), .Y(n2087) );
  INVXLTH U1756 ( .A(n1422), .Y(n2088) );
  INVXLTH U1757 ( .A(n2088), .Y(n2089) );
  INVXLTH U1758 ( .A(n2088), .Y(n2090) );
  INVXLTH U1759 ( .A(n1432), .Y(n2091) );
  INVXLTH U1760 ( .A(n2091), .Y(n2092) );
  INVXLTH U1761 ( .A(n2091), .Y(n2093) );
  INVXLTH U1762 ( .A(n1444), .Y(n2094) );
  INVXLTH U1763 ( .A(n2094), .Y(n2095) );
  INVXLTH U1764 ( .A(n2094), .Y(n2096) );
  INVXLTH U1765 ( .A(n1450), .Y(n2097) );
  INVXLTH U1766 ( .A(n2097), .Y(n2098) );
  INVXLTH U1767 ( .A(n2097), .Y(n2099) );
  INVXLTH U1768 ( .A(n1381), .Y(n2100) );
  INVXLTH U1769 ( .A(n2100), .Y(n2101) );
  INVXLTH U1770 ( .A(n2100), .Y(n2102) );
  INVXLTH U1771 ( .A(n1384), .Y(n2103) );
  INVXLTH U1772 ( .A(n2103), .Y(n2104) );
  INVXLTH U1773 ( .A(n2103), .Y(n2105) );
  INVXLTH U1774 ( .A(n1406), .Y(n2106) );
  INVXLTH U1775 ( .A(n2106), .Y(n2107) );
  INVXLTH U1776 ( .A(n2106), .Y(n2108) );
  INVXLTH U1777 ( .A(n1410), .Y(n2109) );
  INVXLTH U1778 ( .A(n2109), .Y(n2110) );
  INVXLTH U1779 ( .A(n2109), .Y(n2111) );
  INVXLTH U1780 ( .A(n1436), .Y(n2112) );
  INVXLTH U1781 ( .A(n2112), .Y(n2113) );
  INVXLTH U1782 ( .A(n2112), .Y(n2114) );
  INVXLTH U1783 ( .A(n1423), .Y(n2115) );
  INVXLTH U1784 ( .A(n2115), .Y(n2116) );
  INVXLTH U1785 ( .A(n2115), .Y(n2117) );
  INVXLTH U1786 ( .A(n1417), .Y(n2118) );
  INVXLTH U1787 ( .A(n2118), .Y(n2119) );
  INVXLTH U1788 ( .A(n2118), .Y(n2120) );
  INVXLTH U1789 ( .A(n1440), .Y(n2121) );
  INVXLTH U1790 ( .A(n2121), .Y(n2122) );
  INVXLTH U1791 ( .A(n2121), .Y(n2123) );
  INVXLTH U1792 ( .A(n1403), .Y(n2124) );
  INVXLTH U1793 ( .A(n2124), .Y(n2125) );
  INVXLTH U1794 ( .A(n2124), .Y(n2126) );
  INVXLTH U1795 ( .A(n1369), .Y(n2127) );
  INVXLTH U1796 ( .A(n2127), .Y(n2128) );
  INVXLTH U1797 ( .A(n2127), .Y(n2129) );
  INVXLTH U1798 ( .A(n1386), .Y(n2130) );
  INVXLTH U1799 ( .A(n2130), .Y(n2131) );
  INVXLTH U1800 ( .A(n2130), .Y(n2132) );
  INVXLTH U1801 ( .A(n1397), .Y(n2133) );
  INVXLTH U1802 ( .A(n2133), .Y(n2134) );
  INVXLTH U1803 ( .A(n2133), .Y(n2135) );
  INVXLTH U1804 ( .A(n1373), .Y(n2136) );
  INVXLTH U1805 ( .A(n2136), .Y(n2137) );
  INVXLTH U1806 ( .A(n2136), .Y(n2138) );
  INVXLTH U1807 ( .A(n1452), .Y(n2139) );
  INVXLTH U1808 ( .A(n2139), .Y(n2140) );
  INVXLTH U1809 ( .A(n2139), .Y(n2141) );
  INVXLTH U1810 ( .A(n1389), .Y(n2142) );
  INVXLTH U1811 ( .A(n2142), .Y(n2143) );
  INVXLTH U1812 ( .A(n2142), .Y(n2144) );
  INVXLTH U1813 ( .A(n1459), .Y(n2145) );
  INVXLTH U1814 ( .A(n2145), .Y(n2146) );
  INVXLTH U1815 ( .A(n2145), .Y(n2147) );
  INVXLTH U1816 ( .A(n1416), .Y(n2148) );
  INVXLTH U1817 ( .A(n2148), .Y(n2149) );
  INVXLTH U1818 ( .A(n2148), .Y(n2150) );
  INVXLTH U1819 ( .A(n1457), .Y(n2151) );
  INVXLTH U1820 ( .A(n2151), .Y(n2152) );
  INVXLTH U1821 ( .A(n2151), .Y(n2153) );
  INVXLTH U1822 ( .A(n1434), .Y(n2154) );
  INVXLTH U1823 ( .A(n2154), .Y(n2155) );
  INVXLTH U1824 ( .A(n2154), .Y(n2156) );
  INVXLTH U1825 ( .A(n1442), .Y(n2157) );
  INVXLTH U1826 ( .A(n2157), .Y(n2158) );
  INVXLTH U1827 ( .A(n2157), .Y(n2159) );
  INVXLTH U1828 ( .A(n1428), .Y(n2160) );
  INVXLTH U1829 ( .A(n2160), .Y(n2161) );
  INVXLTH U1830 ( .A(n2160), .Y(n2162) );
  INVXLTH U1831 ( .A(n1429), .Y(n2163) );
  INVXLTH U1832 ( .A(n2163), .Y(n2164) );
  INVXLTH U1833 ( .A(n2163), .Y(n2165) );
  INVXLTH U1834 ( .A(n1447), .Y(n2166) );
  INVXLTH U1835 ( .A(n2166), .Y(n2167) );
  INVXLTH U1836 ( .A(n2166), .Y(n2168) );
  INVXLTH U1837 ( .A(n1448), .Y(n2169) );
  INVXLTH U1838 ( .A(n2169), .Y(n2170) );
  INVXLTH U1839 ( .A(n2169), .Y(n2171) );
  INVXLTH U1840 ( .A(n1445), .Y(n2172) );
  INVXLTH U1841 ( .A(n2172), .Y(n2173) );
  INVXLTH U1842 ( .A(n2172), .Y(n2174) );
  INVXLTH U1843 ( .A(n1446), .Y(n2175) );
  INVXLTH U1844 ( .A(n2175), .Y(n2176) );
  INVXLTH U1845 ( .A(n2175), .Y(n2177) );
  INVXLTH U1846 ( .A(n1415), .Y(n2178) );
  INVXLTH U1847 ( .A(n2178), .Y(n2179) );
  INVXLTH U1848 ( .A(n2178), .Y(n2180) );
  INVXLTH U1849 ( .A(n1421), .Y(n2181) );
  INVXLTH U1850 ( .A(n2181), .Y(n2182) );
  INVXLTH U1851 ( .A(n2181), .Y(n2183) );
  INVXLTH U1852 ( .A(n1439), .Y(n2184) );
  INVXLTH U1853 ( .A(n2184), .Y(n2185) );
  INVXLTH U1854 ( .A(n2184), .Y(n2186) );
  INVXLTH U1855 ( .A(n1426), .Y(n2187) );
  INVXLTH U1856 ( .A(n2187), .Y(n2188) );
  INVXLTH U1857 ( .A(n2187), .Y(n2189) );
  INVXLTH U1858 ( .A(n1449), .Y(n2190) );
  INVXLTH U1859 ( .A(n2190), .Y(n2191) );
  INVXLTH U1860 ( .A(n2190), .Y(n2192) );
  INVXLTH U1861 ( .A(n1431), .Y(n2193) );
  INVXLTH U1862 ( .A(n2193), .Y(n2194) );
  INVXLTH U1863 ( .A(n2193), .Y(n2195) );
  INVXLTH U1864 ( .A(n1427), .Y(n2196) );
  INVXLTH U1865 ( .A(n2196), .Y(n2197) );
  INVXLTH U1866 ( .A(n2196), .Y(n2198) );
  INVXLTH U1867 ( .A(n1438), .Y(n2199) );
  INVXLTH U1868 ( .A(n2199), .Y(n2200) );
  INVXLTH U1869 ( .A(n2199), .Y(n2201) );
  INVXLTH U1870 ( .A(n1435), .Y(n2202) );
  INVXLTH U1871 ( .A(n2202), .Y(n2203) );
  INVXLTH U1872 ( .A(n2202), .Y(n2204) );
  INVXLTH U1873 ( .A(n1409), .Y(n2205) );
  INVXLTH U1874 ( .A(n2205), .Y(n2206) );
  INVXLTH U1875 ( .A(n2205), .Y(n2207) );
  INVXLTH U1876 ( .A(n1430), .Y(n2208) );
  INVXLTH U1877 ( .A(n2208), .Y(n2209) );
  INVXLTH U1878 ( .A(n2208), .Y(n2210) );
  INVXLTH U1879 ( .A(n1412), .Y(n2211) );
  INVXLTH U1880 ( .A(n2211), .Y(n2212) );
  INVXLTH U1881 ( .A(n2211), .Y(n2213) );
  INVXLTH U1882 ( .A(n1443), .Y(n2214) );
  INVXLTH U1883 ( .A(n2214), .Y(n2215) );
  INVXLTH U1884 ( .A(n2214), .Y(n2216) );
  INVXLTH U1885 ( .A(n1413), .Y(n2217) );
  INVXLTH U1886 ( .A(n2217), .Y(n2218) );
  INVXLTH U1887 ( .A(n2217), .Y(n2219) );
  INVXLTH U1888 ( .A(n1405), .Y(n2220) );
  INVXLTH U1889 ( .A(n2220), .Y(n2221) );
  INVXLTH U1890 ( .A(n2220), .Y(n2222) );
  INVXLTH U1891 ( .A(n1453), .Y(n2223) );
  INVXLTH U1892 ( .A(n2223), .Y(n2224) );
  INVXLTH U1893 ( .A(n2223), .Y(n2225) );
  INVXLTH U1894 ( .A(n1394), .Y(n2226) );
  INVXLTH U1895 ( .A(n2226), .Y(n2227) );
  INVXLTH U1896 ( .A(n2226), .Y(n2228) );
  INVXLTH U1897 ( .A(n1375), .Y(n2229) );
  INVXLTH U1898 ( .A(n2229), .Y(n2230) );
  INVXLTH U1899 ( .A(n2229), .Y(n2231) );
  INVXLTH U1900 ( .A(n1376), .Y(n2232) );
  INVXLTH U1901 ( .A(n2232), .Y(n2233) );
  INVXLTH U1902 ( .A(n2232), .Y(n2234) );
  INVXLTH U1903 ( .A(n1400), .Y(n2235) );
  INVXLTH U1904 ( .A(n2235), .Y(n2236) );
  INVXLTH U1905 ( .A(n2235), .Y(n2237) );
  INVXLTH U1906 ( .A(n1402), .Y(n2238) );
  INVXLTH U1907 ( .A(n2238), .Y(n2239) );
  INVXLTH U1908 ( .A(n2238), .Y(n2240) );
  INVXLTH U1909 ( .A(n1372), .Y(n2241) );
  INVXLTH U1910 ( .A(n2241), .Y(n2242) );
  INVXLTH U1911 ( .A(n2241), .Y(n2243) );
  INVXLTH U1912 ( .A(n1388), .Y(n2244) );
  INVXLTH U1913 ( .A(n2244), .Y(n2245) );
  INVXLTH U1914 ( .A(n2244), .Y(n2246) );
  INVXLTH U1915 ( .A(n1278), .Y(n2247) );
  INVXLTH U1916 ( .A(n2247), .Y(n2248) );
  INVXLTH U1917 ( .A(n2247), .Y(n2249) );
  INVXLTH U1918 ( .A(n1321), .Y(n2250) );
  INVXLTH U1919 ( .A(n2250), .Y(n2251) );
  INVXLTH U1920 ( .A(n2250), .Y(n2252) );
  INVXLTH U1921 ( .A(n1229), .Y(n2253) );
  INVXLTH U1922 ( .A(n2253), .Y(n2254) );
  INVXLTH U1923 ( .A(n2253), .Y(n2255) );
  INVXLTH U1924 ( .A(n1322), .Y(n2256) );
  INVXLTH U1925 ( .A(n2256), .Y(n2257) );
  INVXLTH U1926 ( .A(n2256), .Y(n2258) );
  INVXLTH U1927 ( .A(n1236), .Y(n2259) );
  INVXLTH U1928 ( .A(n2259), .Y(n2260) );
  INVXLTH U1929 ( .A(n2259), .Y(n2261) );
  DLY1X1TH U1930 ( .A(out47[2]), .Y(n2262) );
  DLY1X1TH U1931 ( .A(out0[4]), .Y(n2263) );
endmodule


module awgn_gen_test_1 ( out1, out2, out3, out4, out5, out6, out7, out8, out9, 
        out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, 
        out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, 
        out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, 
        out40, out41, out42, out43, out44, out45, out46, out47, out48, count1, 
        count2, ex_clk, reset, db, codeword, reset_lfsr, data_sel, data_in, 
        test_si, test_so, test_se );
  output [4:0] out1;
  output [4:0] out2;
  output [4:0] out3;
  output [4:0] out4;
  output [4:0] out5;
  output [4:0] out6;
  output [4:0] out7;
  output [4:0] out8;
  output [4:0] out9;
  output [4:0] out10;
  output [4:0] out11;
  output [4:0] out12;
  output [4:0] out13;
  output [4:0] out14;
  output [4:0] out15;
  output [4:0] out16;
  output [4:0] out17;
  output [4:0] out18;
  output [4:0] out19;
  output [4:0] out20;
  output [4:0] out21;
  output [4:0] out22;
  output [4:0] out23;
  output [4:0] out24;
  output [4:0] out25;
  output [4:0] out26;
  output [4:0] out27;
  output [4:0] out28;
  output [4:0] out29;
  output [4:0] out30;
  output [4:0] out31;
  output [4:0] out32;
  output [4:0] out33;
  output [4:0] out34;
  output [4:0] out35;
  output [4:0] out36;
  output [4:0] out37;
  output [4:0] out38;
  output [4:0] out39;
  output [4:0] out40;
  output [4:0] out41;
  output [4:0] out42;
  output [4:0] out43;
  output [4:0] out44;
  output [4:0] out45;
  output [4:0] out46;
  output [4:0] out47;
  output [4:0] out48;
  output [9:0] count2;
  input [2:0] db;
  input [4:0] data_in;
  input ex_clk, reset, codeword, reset_lfsr, data_sel, test_si, test_se;
  output count1, test_so;
  wire   n3, n4, n8, n9, n10;
  wire   [4:0] qu_llr;
  wire   [4:0] qu_llrr;

  awgn_test_1 awgn_1 ( .clk(ex_clk), .reset(n3), .db(db), .qu_llr(qu_llr), 
        .codeword(codeword), .test_si(out48[4]), .test_so(test_so), .test_se(
        n9) );
  data_mux data_mux_1 ( .out(qu_llrr), .in1(data_in), .in2(qu_llr), .sel(
        data_sel) );
  SIPO_test_1 SIPO_1 ( .out0(out1), .out1(out2), .out2(out3), .out3(out4), 
        .out4(out5), .out5(out6), .out6(out7), .out7(out8), .out8(out9), 
        .out9(out10), .out10(out11), .out11(out12), .out12(out13), .out13(
        out14), .out14(out15), .out15(out16), .out16(out17), .out17(out18), 
        .out18(out19), .out19(out20), .out20(out21), .out21(out22), .out22(
        out23), .out23(out24), .out24(out25), .out25(out26), .out26(out27), 
        .out27(out28), .out28(out29), .out29(out30), .out30(out31), .out31(
        out32), .out32(out33), .out33(out34), .out34(out35), .out35(out36), 
        .out36(out37), .out37(out38), .out38(out39), .out39(out40), .out40(
        out41), .out41(out42), .out42(out43), .out43(out44), .out44(out45), 
        .out45(out46), .out46(out47), .out47(out48), .count1(count1), .count2(
        count2), .in(qu_llrr), .reset(n4), .clk(ex_clk), .test_si(test_si), 
        .test_se(n10) );
  CLKBUFX1TH U1 ( .A(reset), .Y(n4) );
  CLKBUFX1TH U2 ( .A(reset_lfsr), .Y(n3) );
  INVXLTH U3 ( .A(test_se), .Y(n8) );
  INVXLTH U4 ( .A(n8), .Y(n9) );
  INVXLTH U5 ( .A(n8), .Y(n10) );
endmodule


module full_ldpc_decoder_test_1 ( error_codeword, error, hd_end, in_clk, 
        iteration_start, iteration_end, out_hd, db, codeword, sel, ex_clk, rst, 
        reset_lfsr, TM, data_sel, data_in, test_si, test_so, test_se );
  output [9:0] error_codeword;
  output [9:0] error;
  input [2:0] db;
  input [1:0] sel;
  input [4:0] data_in;
  input codeword, ex_clk, rst, reset_lfsr, TM, data_sel, test_si, test_se;
  output hd_end, in_clk, iteration_start, iteration_end, out_hd, test_so;
  wire   intt_clk, int_clk, out1, out2, out3, out4, out5, out6, out7, out8,
         out9, out10, out11, out12, out13, out14, out15, out16, out17, out18,
         out19, out20, out21, out22, out23, out24, out25, out26, out27, out28,
         out29, out30, out31, out32, out33, out34, out35, out36, out37, out38,
         out39, out40, out41, out42, out43, out44, out45, out46, out47, out48,
         n22, n15, n16, n17, n18, n19, n21, n25, n26, n27, n30;
  wire   [4:0] qu_llr1;
  wire   [4:0] qu_llr2;
  wire   [4:0] qu_llr3;
  wire   [4:0] qu_llr4;
  wire   [4:0] qu_llr5;
  wire   [4:0] qu_llr6;
  wire   [4:0] qu_llr7;
  wire   [4:0] qu_llr8;
  wire   [4:0] qu_llr9;
  wire   [4:0] qu_llr10;
  wire   [4:0] qu_llr11;
  wire   [4:0] qu_llr12;
  wire   [4:0] qu_llr13;
  wire   [4:0] qu_llr14;
  wire   [4:0] qu_llr15;
  wire   [4:0] qu_llr16;
  wire   [4:0] qu_llr17;
  wire   [4:0] qu_llr18;
  wire   [4:0] qu_llr19;
  wire   [4:0] qu_llr20;
  wire   [4:0] qu_llr21;
  wire   [4:0] qu_llr22;
  wire   [4:0] qu_llr23;
  wire   [4:0] qu_llr24;
  wire   [4:0] qu_llr25;
  wire   [4:0] qu_llr26;
  wire   [4:0] qu_llr27;
  wire   [4:0] qu_llr28;
  wire   [4:0] qu_llr29;
  wire   [4:0] qu_llr30;
  wire   [4:0] qu_llr31;
  wire   [4:0] qu_llr32;
  wire   [4:0] qu_llr33;
  wire   [4:0] qu_llr34;
  wire   [4:0] qu_llr35;
  wire   [4:0] qu_llr36;
  wire   [4:0] qu_llr37;
  wire   [4:0] qu_llr38;
  wire   [4:0] qu_llr39;
  wire   [4:0] qu_llr40;
  wire   [4:0] qu_llr41;
  wire   [4:0] qu_llr42;
  wire   [4:0] qu_llr43;
  wire   [4:0] qu_llr44;
  wire   [4:0] qu_llr45;
  wire   [4:0] qu_llr46;
  wire   [4:0] qu_llr47;
  wire   [4:0] qu_llr48;

  TLATNTSCAX6 TLATNTSCAX6_1 ( .E(iteration_start), .SE(TM), .CK(ex_clk), .ECK(
        int_clk) );
  fmod4_test_1 fmod4_1 ( .out(intt_clk), .clk(ex_clk), .rst(n17), .test_si(
        hd_end), .test_so(n25), .test_se(test_se) );
  mux_top mux_top_1 ( .out(in_clk), .in1(ex_clk), .in2(intt_clk), .sel(TM) );
  awgn_gen_test_1 awrn_gen_1 ( .out1(qu_llr1), .out2(qu_llr2), .out3(qu_llr3), 
        .out4(qu_llr4), .out5(qu_llr5), .out6(qu_llr6), .out7(qu_llr7), .out8(
        qu_llr8), .out9(qu_llr9), .out10(qu_llr10), .out11(qu_llr11), .out12(
        qu_llr12), .out13(qu_llr13), .out14(qu_llr14), .out15(qu_llr15), 
        .out16(qu_llr16), .out17(qu_llr17), .out18(qu_llr18), .out19(qu_llr19), 
        .out20(qu_llr20), .out21(qu_llr21), .out22(qu_llr22), .out23(qu_llr23), 
        .out24(qu_llr24), .out25(qu_llr25), .out26(qu_llr26), .out27(qu_llr27), 
        .out28(qu_llr28), .out29(qu_llr29), .out30(qu_llr30), .out31(qu_llr31), 
        .out32(qu_llr32), .out33(qu_llr33), .out34(qu_llr34), .out35(qu_llr35), 
        .out36(qu_llr36), .out37(qu_llr37), .out38(qu_llr38), .out39(qu_llr39), 
        .out40(qu_llr40), .out41(qu_llr41), .out42(qu_llr42), .out43(qu_llr43), 
        .out44(qu_llr44), .out45(qu_llr45), .out46(qu_llr46), .out47(qu_llr47), 
        .out48(qu_llr48), .count1(iteration_start), .count2(error_codeword), 
        .ex_clk(in_clk), .reset(n18), .db(db), .codeword(codeword), 
        .reset_lfsr(reset_lfsr), .data_sel(data_sel), .data_in(data_in), 
        .test_si(test_si), .test_so(n27), .test_se(test_se) );
  counter_test_1 counter_1 ( .out1(n22), .sel(sel), .clk(int_clk), .rst(rst), 
        .test_si(n27), .test_so(n26), .test_se(n30) );
  counter_PISO_test_1 counter_PISO_1 ( .error(error), .hd_end(hd_end), .in1(
        out1), .in2(out2), .in3(out3), .in4(out4), .in5(out5), .in6(out6), 
        .in7(out7), .in8(out8), .in9(out9), .in10(out10), .in11(out11), .in12(
        out12), .in13(out13), .in14(out14), .in15(out15), .in16(out16), .in17(
        out17), .in18(out18), .in19(out19), .in20(out20), .in21(out21), .in22(
        out22), .in23(out23), .in24(out24), .in25(out25), .in26(out26), .in27(
        out27), .in28(out28), .in29(out29), .in30(out30), .in31(out31), .in32(
        out32), .in33(out33), .in34(out34), .in35(out35), .in36(out36), .in37(
        out37), .in38(out38), .in39(out39), .in40(out40), .in41(out41), .in42(
        out42), .in43(out43), .in44(out44), .in45(out45), .in46(out46), .in47(
        out47), .in48(out48), .rst(n16), .ex_clk(int_clk), .w3(iteration_end), 
        .test_si(n26), .test_se(test_se) );
  iteration_test_1 iter1 ( .h1(out1), .h2(out2), .h3(out3), .h4(out4), .h5(
        out5), .h6(out6), .h7(out7), .h8(out8), .h9(out9), .h10(out10), .h11(
        out11), .h12(out12), .h13(out13), .h14(out14), .h15(out15), .h16(out16), .h17(out17), .h18(out18), .h19(out19), .h20(out20), .h21(out21), .h22(out22), 
        .h23(out23), .h24(out24), .h25(out25), .h26(out26), .h27(out27), .h28(
        out28), .h29(out29), .h30(out30), .h31(out31), .h32(out32), .h33(out33), .h34(out34), .h35(out35), .h36(out36), .h37(out37), .h38(out38), .h39(out39), 
        .h40(out40), .h41(out41), .h42(out42), .h43(out43), .h44(out44), .h45(
        out45), .h46(out46), .h47(out47), .h48(out48), .clk(int_clk), .rst(n18), .i1(qu_llr1), .i2(qu_llr2), .i3(qu_llr3), .i4(qu_llr4), .i5(qu_llr5), .i6(
        qu_llr6), .i7(qu_llr7), .i8(qu_llr8), .i9(qu_llr9), .i10(qu_llr10), 
        .i11(qu_llr11), .i12(qu_llr12), .i13(qu_llr13), .i14(qu_llr14), .i15(
        qu_llr15), .i16(qu_llr16), .i17(qu_llr17), .i18(qu_llr18), .i19(
        qu_llr19), .i20(qu_llr20), .i21(qu_llr21), .i22(qu_llr22), .i23(
        qu_llr23), .i24(qu_llr24), .i25(qu_llr25), .i26(qu_llr26), .i27(
        qu_llr27), .i28(qu_llr28), .i29(qu_llr29), .i30(qu_llr30), .i31(
        qu_llr31), .i32(qu_llr32), .i33(qu_llr33), .i34(qu_llr34), .i35(
        qu_llr35), .i36(qu_llr36), .i37(qu_llr37), .i38(qu_llr38), .i39(
        qu_llr39), .i40(qu_llr40), .i41(qu_llr41), .i42(qu_llr42), .i43(
        qu_llr43), .i44(qu_llr44), .i45(qu_llr45), .i46(qu_llr46), .i47(
        qu_llr47), .i48(qu_llr48), .test_si(n25), .test_so(test_so), .test_se(
        test_se) );
  INVX2TH U2 ( .A(1'b1), .Y(out_hd) );
  INVXLTH U4 ( .A(n18), .Y(n15) );
  CLKINVX1TH U5 ( .A(n19), .Y(n18) );
  INVXLTH U6 ( .A(n15), .Y(n16) );
  INVXLTH U7 ( .A(n15), .Y(n17) );
  INVXLTH U8 ( .A(n21), .Y(iteration_end) );
  INVXLTH U9 ( .A(n22), .Y(n21) );
  INVXLTH U10 ( .A(rst), .Y(n19) );
  DLY1X1TH U1 ( .A(test_se), .Y(n30) );
endmodule


module CHIP ( error_codeword, error, hd_end, in_clk, iteration_start, 
        iteration_end, out_hd, db, codeword, sel, ex_clk, rst, reset_lfsr, TM, 
        si, so, se, data_sel, data_in );
  output [9:0] error_codeword;
  output [9:0] error;
  input [2:0] db;
  input [1:0] sel;
  input [4:0] data_in;
  input codeword, ex_clk, rst, reset_lfsr, TM, si, se, data_sel;
  output hd_end, in_clk, iteration_start, iteration_end, out_hd, so;
  wire   i_hd_end, i_in_clk, i_iteration_start, i_iteration_end, i_codeword,
         i_ex_clk, i_rst, i_reset_lfsr, i_TM, i_data_sel, n3, n4, n5, n6;
  wire   [9:0] i_error_codeword;
  wire   [9:0] i_error;
  wire   [2:0] i_db;
  wire   [1:0] i_sel;
  wire   [4:0] i_data_in;

  PDO16CDG_33 opad_ERROR_CODEWORD0 ( .I(i_error_codeword[0]), .PAD(
        error_codeword[0]) );
  PDO16CDG_33 opad_ERROR_CODEWORD1 ( .I(i_error_codeword[1]), .PAD(
        error_codeword[1]) );
  PDO16CDG_33 opad_ERROR_CODEWORD2 ( .I(i_error_codeword[2]), .PAD(
        error_codeword[2]) );
  PDO16CDG_33 opad_ERROR_CODEWORD3 ( .I(i_error_codeword[3]), .PAD(
        error_codeword[3]) );
  PDO16CDG_33 opad_ERROR_CODEWORD4 ( .I(i_error_codeword[4]), .PAD(
        error_codeword[4]) );
  PDO16CDG_33 opad_ERROR_CODEWORD5 ( .I(i_error_codeword[5]), .PAD(
        error_codeword[5]) );
  PDO16CDG_33 opad_ERROR_CODEWORD6 ( .I(i_error_codeword[6]), .PAD(
        error_codeword[6]) );
  PDO16CDG_33 opad_ERROR_CODEWORD7 ( .I(i_error_codeword[7]), .PAD(
        error_codeword[7]) );
  PDO16CDG_33 opad_ERROR_CODEWORD8 ( .I(i_error_codeword[8]), .PAD(
        error_codeword[8]) );
  PDO16CDG_33 opad_ERROR_CODEWORD9 ( .I(i_error_codeword[9]), .PAD(
        error_codeword[9]) );
  PDO16CDG_33 opad_ERROR0 ( .I(i_error[0]), .PAD(error[0]) );
  PDO16CDG_33 opad_ERROR1 ( .I(i_error[1]), .PAD(error[1]) );
  PDO16CDG_33 opad_ERROR2 ( .I(i_error[2]), .PAD(error[2]) );
  PDO16CDG_33 opad_ERROR3 ( .I(i_error[3]), .PAD(error[3]) );
  PDO16CDG_33 opad_ERROR4 ( .I(i_error[4]), .PAD(error[4]) );
  PDO16CDG_33 opad_ERROR5 ( .I(i_error[5]), .PAD(error[5]) );
  PDO16CDG_33 opad_ERROR6 ( .I(i_error[6]), .PAD(error[6]) );
  PDO16CDG_33 opad_ERROR7 ( .I(i_error[7]), .PAD(error[7]) );
  PDO16CDG_33 opad_ERROR8 ( .I(i_error[8]), .PAD(error[8]) );
  PDO16CDG_33 opad_ERROR9 ( .I(i_error[9]), .PAD(error[9]) );
  PDO16CDG_33 opad_HD_END ( .I(i_hd_end), .PAD(hd_end) );
  PDO16CDG_33 opad_IN_CLK ( .I(i_in_clk), .PAD(in_clk) );
  PDO16CDG_33 opad_ITERATION_START ( .I(i_iteration_start), .PAD(
        iteration_start) );
  PDO16CDG_33 opad_ITERATION_END ( .I(n3), .PAD(iteration_end) );
  PDO16CDG_33 opad_OUT_HD ( .I(1'b0), .PAD(out_hd) );
  PDO16CDG_33 opad_SO ( .I(n5), .PAD(so) );
  PDIDGZ_33 ipad_DB0 ( .PAD(db[0]), .C(i_db[0]) );
  PDIDGZ_33 ipad_DB1 ( .PAD(db[1]), .C(i_db[1]) );
  PDIDGZ_33 ipad_DB2 ( .PAD(db[2]), .C(i_db[2]) );
  PDIDGZ_33 ipad_CODEWORD ( .PAD(codeword), .C(i_codeword) );
  PDIDGZ_33 ipad_SEL0 ( .PAD(sel[0]), .C(i_sel[0]) );
  PDIDGZ_33 ipad_SEL1 ( .PAD(sel[1]), .C(i_sel[1]) );
  PDIDGZ_33 ipad_EX_CLK ( .PAD(ex_clk), .C(i_ex_clk) );
  PDIDGZ_33 ipad_RST ( .PAD(rst), .C(i_rst) );
  PDIDGZ_33 ipad_RESET_LFSR ( .PAD(reset_lfsr), .C(i_reset_lfsr) );
  PDIDGZ_33 ipad_TM ( .PAD(TM), .C(i_TM) );
  PDIDGZ_33 ipad_SI ( .PAD(si), .C(n6) );
  PDIDGZ_33 ipad_SE ( .PAD(se), .C(n4) );
  PDIDGZ_33 ipad_DATA_IN0 ( .PAD(data_in[0]), .C(i_data_in[0]) );
  PDIDGZ_33 ipad_DATA_IN1 ( .PAD(data_in[1]), .C(i_data_in[1]) );
  PDIDGZ_33 ipad_DATA_IN2 ( .PAD(data_in[2]), .C(i_data_in[2]) );
  PDIDGZ_33 ipad_DATA_IN3 ( .PAD(data_in[3]), .C(i_data_in[3]) );
  PDIDGZ_33 ipad_DATA_IN4 ( .PAD(data_in[4]), .C(i_data_in[4]) );
  PDIDGZ_33 ipad_DATA_SEL ( .PAD(data_sel), .C(i_data_sel) );
  full_ldpc_decoder_test_1 full_ldpc_decoder_1 ( .error_codeword(
        i_error_codeword), .error(i_error), .hd_end(i_hd_end), .in_clk(
        i_in_clk), .iteration_start(i_iteration_start), .iteration_end(
        i_iteration_end), .db(i_db), .codeword(i_codeword), .sel(i_sel), 
        .ex_clk(i_ex_clk), .rst(i_rst), .reset_lfsr(i_reset_lfsr), .TM(i_TM), 
        .data_sel(i_data_sel), .data_in(i_data_in), .test_si(n6), .test_so(n5), 
        .test_se(n4) );
  CLKBUFX2TH U1 ( .A(i_iteration_end), .Y(n3) );
endmodule

